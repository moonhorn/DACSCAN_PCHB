//
// bench2vlog.py
//   options: -l nangate --clk CK --si test_si --so test_so --se test_se
//
module s38417 (CK,  g51, g563, g1249, g1943, g2637, g3212, g3213, g3214, g3215, g3216, g3217, g3218, g3219, g3220, g3221, g3222, g3223, g3224, g3225, g3226, g3227, g3228, g3229, g3230, g3231, g3232, g3233, g3234, g3993, g4088, g4090, g4200, g4321, g4323, g4450, g4590, g5388, g5437, g5472, g5511, g5549, g5555, g5595, g5612, g5629, g5637, g5648, g5657, g5686, g5695, g5738, g5747, g5796, g6225, g6231, g6313, g6368, g6442, g6447, g6485, g6518, g6573, g6642, g6677, g6712, g6750, g6782, g6837, g6895, g6911, g6944, g6979, g7014, g7052, g7084, g7161, g7194, g7229, g7264, g7302, g7334, g7357, g7390, g7425, g7487, g7519, g7909, g7956, g7961, g8007, g8012, g8021, g8023, g8030, g8082, g8087, g8096, g8106, g8167, g8175, g8249, g8251, g8258, g8259, g8260, g8261, g8262, g8263, g8264, g8265, g8266, g8267, g8268, g8269, g8270, g8271, g8272, g8273, g8274, g8275, g16297, g16355, g16399, g16437, g16496, g24734, g25420, g25435, g25442, g25489, g26104, g26135, g26149, g27380);

input g51 ;
input g563 ;
input g1249 ;
input g1943 ;
input g2637 ;
input g3212 ;
input g3213 ;
input g3214 ;
input g3215 ;
input g3216 ;
input g3217 ;
input g3218 ;
input g3219 ;
input g3220 ;
input g3221 ;
input g3222 ;
input g3223 ;
input g3224 ;
input g3225 ;
input g3226 ;
input g3227 ;
input g3228 ;
input g3229 ;
input g3230 ;
input g3231 ;
input g3232 ;
input g3233 ;
input g3234 ;
input CK ;

output g3993 ;
output g4088 ;
output g4090 ;
output g4200 ;
output g4321 ;
output g4323 ;
output g4450 ;
output g4590 ;
output g5388 ;
output g5437 ;
output g5472 ;
output g5511 ;
output g5549 ;
output g5555 ;
output g5595 ;
output g5612 ;
output g5629 ;
output g5637 ;
output g5648 ;
output g5657 ;
output g5686 ;
output g5695 ;
output g5738 ;
output g5747 ;
output g5796 ;
output g6225 ;
output g6231 ;
output g6313 ;
output g6368 ;
output g6442 ;
output g6447 ;
output g6485 ;
output g6518 ;
output g6573 ;
output g6642 ;
output g6677 ;
output g6712 ;
output g6750 ;
output g6782 ;
output g6837 ;
output g6895 ;
output g6911 ;
output g6944 ;
output g6979 ;
output g7014 ;
output g7052 ;
output g7084 ;
output g7161 ;
output g7194 ;
output g7229 ;
output g7264 ;
output g7302 ;
output g7334 ;
output g7357 ;
output g7390 ;
output g7425 ;
output g7487 ;
output g7519 ;
output g7909 ;
output g7956 ;
output g7961 ;
output g8007 ;
output g8012 ;
output g8021 ;
output g8023 ;
output g8030 ;
output g8082 ;
output g8087 ;
output g8096 ;
output g8106 ;
output g8167 ;
output g8175 ;
output g8249 ;
output g8251 ;
output g8258 ;
output g8259 ;
output g8260 ;
output g8261 ;
output g8262 ;
output g8263 ;
output g8264 ;
output g8265 ;
output g8266 ;
output g8267 ;
output g8268 ;
output g8269 ;
output g8270 ;
output g8271 ;
output g8272 ;
output g8273 ;
output g8274 ;
output g8275 ;
output g16297 ;
output g16355 ;
output g16399 ;
output g16437 ;
output g16496 ;
output g24734 ;
output g25420 ;
output g25435 ;
output g25442 ;
output g25489 ;
output g26104 ;
output g26135 ;
output g26149 ;
output g27380 ;

//startLogic
INV_X32 U_I13089 ( .A(g563), .ZN(I13089) );
INV_X32 U_g562 ( .A(I13089), .ZN(g562) );
INV_X32 U_I13092 ( .A(g1249), .ZN(I13092) );
INV_X32 U_g1248 ( .A(I13092), .ZN(g1248) );
INV_X32 U_I13095 ( .A(g1943), .ZN(I13095) );
INV_X32 U_g1942 ( .A(I13095), .ZN(g1942) );
INV_X32 U_I13098 ( .A(g2637), .ZN(I13098) );
INV_X32 U_g2636 ( .A(I13098), .ZN(g2636) );
INV_X32 U_I13101 ( .A(g1), .ZN(I13101) );
INV_X32 U_g3235 ( .A(I13101), .ZN(g3235) );
INV_X32 U_I13104 ( .A(g2), .ZN(I13104) );
INV_X32 U_g3236 ( .A(I13104), .ZN(g3236) );
INV_X32 U_I13107 ( .A(g5), .ZN(I13107) );
INV_X32 U_g3237 ( .A(I13107), .ZN(g3237) );
INV_X32 U_I13110 ( .A(g8), .ZN(I13110) );
INV_X32 U_g3238 ( .A(I13110), .ZN(g3238) );
INV_X32 U_I13113 ( .A(g11), .ZN(I13113) );
INV_X32 U_g3239 ( .A(I13113), .ZN(g3239) );
INV_X32 U_I13116 ( .A(g14), .ZN(I13116) );
INV_X32 U_g3240 ( .A(I13116), .ZN(g3240) );
INV_X32 U_I13119 ( .A(g17), .ZN(I13119) );
INV_X32 U_g3241 ( .A(I13119), .ZN(g3241) );
INV_X32 U_I13122 ( .A(g20), .ZN(I13122) );
INV_X32 U_g3242 ( .A(I13122), .ZN(g3242) );
INV_X32 U_I13125 ( .A(g23), .ZN(I13125) );
INV_X32 U_g3243 ( .A(I13125), .ZN(g3243) );
INV_X32 U_I13128 ( .A(g26), .ZN(I13128) );
INV_X32 U_g3244 ( .A(I13128), .ZN(g3244) );
INV_X32 U_I13131 ( .A(g27), .ZN(I13131) );
INV_X32 U_g3245 ( .A(I13131), .ZN(g3245) );
INV_X32 U_I13134 ( .A(g30), .ZN(I13134) );
INV_X32 U_g3246 ( .A(I13134), .ZN(g3246) );
INV_X32 U_I13137 ( .A(g33), .ZN(I13137) );
INV_X32 U_g3247 ( .A(I13137), .ZN(g3247) );
INV_X32 U_I13140 ( .A(g36), .ZN(I13140) );
INV_X32 U_g3248 ( .A(I13140), .ZN(g3248) );
INV_X32 U_I13143 ( .A(g39), .ZN(I13143) );
INV_X32 U_g3249 ( .A(I13143), .ZN(g3249) );
INV_X32 U_I13146 ( .A(g42), .ZN(I13146) );
INV_X32 U_g3250 ( .A(I13146), .ZN(g3250) );
INV_X32 U_I13149 ( .A(g45), .ZN(I13149) );
INV_X32 U_g3251 ( .A(I13149), .ZN(g3251) );
INV_X32 U_I13152 ( .A(g48), .ZN(I13152) );
INV_X32 U_g3252 ( .A(I13152), .ZN(g3252) );
INV_X32 U_I13155 ( .A(g51), .ZN(I13155) );
INV_X32 U_g3253 ( .A(I13155), .ZN(g3253) );
INV_X32 U_I13158 ( .A(g165), .ZN(I13158) );
INV_X32 U_g3254 ( .A(I13158), .ZN(g3254) );
INV_X32 U_I13161 ( .A(g308), .ZN(I13161) );
INV_X32 U_g3304 ( .A(I13161), .ZN(g3304) );
INV_X32 U_g3305 ( .A(g305), .ZN(g3305) );
INV_X32 U_I13165 ( .A(g401), .ZN(I13165) );
INV_X32 U_g3306 ( .A(I13165), .ZN(g3306) );
INV_X32 U_g3337 ( .A(g309), .ZN(g3337) );
INV_X32 U_I13169 ( .A(g550), .ZN(I13169) );
INV_X32 U_g3338 ( .A(I13169), .ZN(g3338) );
INV_X32 U_g3365 ( .A(g499), .ZN(g3365) );
INV_X32 U_I13173 ( .A(g629), .ZN(I13173) );
INV_X32 U_g3366 ( .A(I13173), .ZN(g3366) );
INV_X32 U_I13176 ( .A(g630), .ZN(I13176) );
INV_X32 U_g3398 ( .A(I13176), .ZN(g3398) );
INV_X32 U_I13179 ( .A(g853), .ZN(I13179) );
INV_X32 U_g3410 ( .A(I13179), .ZN(g3410) );
INV_X32 U_I13182 ( .A(g995), .ZN(I13182) );
INV_X32 U_g3460 ( .A(I13182), .ZN(g3460) );
INV_X32 U_g3461 ( .A(g992), .ZN(g3461) );
INV_X32 U_I13186 ( .A(g1088), .ZN(I13186) );
INV_X32 U_g3462 ( .A(I13186), .ZN(g3462) );
INV_X32 U_g3493 ( .A(g996), .ZN(g3493) );
INV_X32 U_I13190 ( .A(g1236), .ZN(I13190) );
INV_X32 U_g3494 ( .A(I13190), .ZN(g3494) );
INV_X32 U_g3521 ( .A(g1186), .ZN(g3521) );
INV_X32 U_I13194 ( .A(g1315), .ZN(I13194) );
INV_X32 U_g3522 ( .A(I13194), .ZN(g3522) );
INV_X32 U_I13197 ( .A(g1316), .ZN(I13197) );
INV_X32 U_g3554 ( .A(I13197), .ZN(g3554) );
INV_X32 U_I13200 ( .A(g1547), .ZN(I13200) );
INV_X32 U_g3566 ( .A(I13200), .ZN(g3566) );
INV_X32 U_I13203 ( .A(g1689), .ZN(I13203) );
INV_X32 U_g3616 ( .A(I13203), .ZN(g3616) );
INV_X32 U_g3617 ( .A(g1686), .ZN(g3617) );
INV_X32 U_I13207 ( .A(g1782), .ZN(I13207) );
INV_X32 U_g3618 ( .A(I13207), .ZN(g3618) );
INV_X32 U_g3649 ( .A(g1690), .ZN(g3649) );
INV_X32 U_I13211 ( .A(g1930), .ZN(I13211) );
INV_X32 U_g3650 ( .A(I13211), .ZN(g3650) );
INV_X32 U_g3677 ( .A(g1880), .ZN(g3677) );
INV_X32 U_I13215 ( .A(g2009), .ZN(I13215) );
INV_X32 U_g3678 ( .A(I13215), .ZN(g3678) );
INV_X32 U_I13218 ( .A(g2010), .ZN(I13218) );
INV_X32 U_g3710 ( .A(I13218), .ZN(g3710) );
INV_X32 U_I13221 ( .A(g2241), .ZN(I13221) );
INV_X32 U_g3722 ( .A(I13221), .ZN(g3722) );
INV_X32 U_I13224 ( .A(g2383), .ZN(I13224) );
INV_X32 U_g3772 ( .A(I13224), .ZN(g3772) );
INV_X32 U_g3773 ( .A(g2380), .ZN(g3773) );
INV_X32 U_I13228 ( .A(g2476), .ZN(I13228) );
INV_X32 U_g3774 ( .A(I13228), .ZN(g3774) );
INV_X32 U_g3805 ( .A(g2384), .ZN(g3805) );
INV_X32 U_I13232 ( .A(g2624), .ZN(I13232) );
INV_X32 U_g3806 ( .A(I13232), .ZN(g3806) );
INV_X32 U_g3833 ( .A(g2574), .ZN(g3833) );
INV_X32 U_I13236 ( .A(g2703), .ZN(I13236) );
INV_X32 U_g3834 ( .A(I13236), .ZN(g3834) );
INV_X32 U_I13239 ( .A(g2704), .ZN(I13239) );
INV_X32 U_g3866 ( .A(I13239), .ZN(g3866) );
INV_X32 U_I13242 ( .A(g2879), .ZN(I13242) );
INV_X32 U_g3878 ( .A(I13242), .ZN(g3878) );
INV_X32 U_g3897 ( .A(g2950), .ZN(g3897) );
INV_X32 U_I13246 ( .A(g2987), .ZN(I13246) );
INV_X32 U_g3900 ( .A(I13246), .ZN(g3900) );
INV_X32 U_g3919 ( .A(g3080), .ZN(g3919) );
INV_X32 U_g3922 ( .A(g150), .ZN(g3922) );
INV_X32 U_g3925 ( .A(g155), .ZN(g3925) );
INV_X32 U_g3928 ( .A(g157), .ZN(g3928) );
INV_X32 U_g3931 ( .A(g171), .ZN(g3931) );
INV_X32 U_g3934 ( .A(g176), .ZN(g3934) );
INV_X32 U_g3937 ( .A(g178), .ZN(g3937) );
INV_X32 U_g3940 ( .A(g408), .ZN(g3940) );
INV_X32 U_g3941 ( .A(g455), .ZN(g3941) );
INV_X32 U_g3942 ( .A(g699), .ZN(g3942) );
INV_X32 U_g3945 ( .A(g726), .ZN(g3945) );
INV_X32 U_g3948 ( .A(g835), .ZN(g3948) );
INV_X32 U_g3951 ( .A(g840), .ZN(g3951) );
INV_X32 U_g3954 ( .A(g842), .ZN(g3954) );
INV_X32 U_g3957 ( .A(g856), .ZN(g3957) );
INV_X32 U_g3960 ( .A(g861), .ZN(g3960) );
INV_X32 U_g3963 ( .A(g863), .ZN(g3963) );
INV_X32 U_g3966 ( .A(g1526), .ZN(g3966) );
INV_X32 U_g3969 ( .A(g1531), .ZN(g3969) );
INV_X32 U_g3972 ( .A(g1533), .ZN(g3972) );
INV_X32 U_g3975 ( .A(g1552), .ZN(g3975) );
INV_X32 U_g3978 ( .A(g1554), .ZN(g3978) );
INV_X32 U_g3981 ( .A(g2217), .ZN(g3981) );
INV_X32 U_g3984 ( .A(g2222), .ZN(g3984) );
INV_X32 U_g3987 ( .A(g2224), .ZN(g3987) );
INV_X32 U_g3990 ( .A(g2245), .ZN(g3990) );
INV_X32 U_I13275 ( .A(g2848), .ZN(I13275) );
INV_X32 U_g3993 ( .A(I13275), .ZN(g3993) );
INV_X32 U_g3994 ( .A(g2848), .ZN(g3994) );
INV_X32 U_g3995 ( .A(g3064), .ZN(g3995) );
INV_X32 U_g3996 ( .A(g3073), .ZN(g3996) );
INV_X32 U_g3997 ( .A(g45), .ZN(g3997) );
INV_X32 U_g3998 ( .A(g23), .ZN(g3998) );
INV_X32 U_g3999 ( .A(g3204), .ZN(g3999) );
INV_X32 U_g4000 ( .A(g153), .ZN(g4000) );
INV_X32 U_g4003 ( .A(g158), .ZN(g4003) );
INV_X32 U_g4006 ( .A(g160), .ZN(g4006) );
INV_X32 U_g4009 ( .A(g174), .ZN(g4009) );
INV_X32 U_g4012 ( .A(g179), .ZN(g4012) );
INV_X32 U_g4015 ( .A(g411), .ZN(g4015) );
INV_X32 U_g4016 ( .A(g417), .ZN(g4016) );
INV_X32 U_g4017 ( .A(g427), .ZN(g4017) );
INV_X32 U_g4020 ( .A(g700), .ZN(g4020) );
INV_X32 U_g4023 ( .A(g702), .ZN(g4023) );
INV_X32 U_g4026 ( .A(g727), .ZN(g4026) );
INV_X32 U_g4029 ( .A(g838), .ZN(g4029) );
INV_X32 U_g4032 ( .A(g843), .ZN(g4032) );
INV_X32 U_g4035 ( .A(g845), .ZN(g4035) );
INV_X32 U_g4038 ( .A(g859), .ZN(g4038) );
INV_X32 U_g4041 ( .A(g864), .ZN(g4041) );
INV_X32 U_g4044 ( .A(g866), .ZN(g4044) );
INV_X32 U_g4047 ( .A(g1095), .ZN(g4047) );
INV_X32 U_g4048 ( .A(g1142), .ZN(g4048) );
INV_X32 U_g4049 ( .A(g1385), .ZN(g4049) );
INV_X32 U_g4052 ( .A(g1412), .ZN(g4052) );
INV_X32 U_g4055 ( .A(g1529), .ZN(g4055) );
INV_X32 U_g4058 ( .A(g1534), .ZN(g4058) );
INV_X32 U_g4061 ( .A(g1536), .ZN(g4061) );
INV_X32 U_g4064 ( .A(g1550), .ZN(g4064) );
INV_X32 U_g4067 ( .A(g1555), .ZN(g4067) );
INV_X32 U_g4070 ( .A(g1557), .ZN(g4070) );
INV_X32 U_g4073 ( .A(g2220), .ZN(g4073) );
INV_X32 U_g4076 ( .A(g2225), .ZN(g4076) );
INV_X32 U_g4079 ( .A(g2227), .ZN(g4079) );
INV_X32 U_g4082 ( .A(g2246), .ZN(g4082) );
INV_X32 U_g4085 ( .A(g2248), .ZN(g4085) );
INV_X32 U_I13316 ( .A(g2836), .ZN(I13316) );
INV_X32 U_g4088 ( .A(I13316), .ZN(g4088) );
INV_X32 U_g4089 ( .A(g2836), .ZN(g4089) );
INV_X32 U_I13320 ( .A(g2864), .ZN(I13320) );
INV_X32 U_g4090 ( .A(I13320), .ZN(g4090) );
INV_X32 U_g4091 ( .A(g2864), .ZN(g4091) );
INV_X32 U_g4092 ( .A(g3074), .ZN(g4092) );
INV_X32 U_g4093 ( .A(g33), .ZN(g4093) );
INV_X32 U_g4094 ( .A(g3207), .ZN(g4094) );
INV_X32 U_g4095 ( .A(g130), .ZN(g4095) );
INV_X32 U_g4098 ( .A(g156), .ZN(g4098) );
INV_X32 U_g4101 ( .A(g161), .ZN(g4101) );
INV_X32 U_g4104 ( .A(g163), .ZN(g4104) );
INV_X32 U_g4107 ( .A(g177), .ZN(g4107) );
INV_X32 U_g4110 ( .A(g414), .ZN(g4110) );
INV_X32 U_g4111 ( .A(g420), .ZN(g4111) );
INV_X32 U_g4112 ( .A(g428), .ZN(g4112) );
INV_X32 U_g4115 ( .A(g698), .ZN(g4115) );
INV_X32 U_g4118 ( .A(g703), .ZN(g4118) );
INV_X32 U_g4121 ( .A(g705), .ZN(g4121) );
INV_X32 U_g4124 ( .A(g725), .ZN(g4124) );
INV_X32 U_g4127 ( .A(g841), .ZN(g4127) );
INV_X32 U_g4130 ( .A(g846), .ZN(g4130) );
INV_X32 U_g4133 ( .A(g848), .ZN(g4133) );
INV_X32 U_g4136 ( .A(g862), .ZN(g4136) );
INV_X32 U_g4139 ( .A(g867), .ZN(g4139) );
INV_X32 U_g4142 ( .A(g1098), .ZN(g4142) );
INV_X32 U_g4143 ( .A(g1104), .ZN(g4143) );
INV_X32 U_g4144 ( .A(g1114), .ZN(g4144) );
INV_X32 U_g4147 ( .A(g1386), .ZN(g4147) );
INV_X32 U_g4150 ( .A(g1388), .ZN(g4150) );
INV_X32 U_g4153 ( .A(g1413), .ZN(g4153) );
INV_X32 U_g4156 ( .A(g1532), .ZN(g4156) );
INV_X32 U_g4159 ( .A(g1537), .ZN(g4159) );
INV_X32 U_g4162 ( .A(g1539), .ZN(g4162) );
INV_X32 U_g4165 ( .A(g1553), .ZN(g4165) );
INV_X32 U_g4168 ( .A(g1558), .ZN(g4168) );
INV_X32 U_g4171 ( .A(g1560), .ZN(g4171) );
INV_X32 U_g4174 ( .A(g1789), .ZN(g4174) );
INV_X32 U_g4175 ( .A(g1836), .ZN(g4175) );
INV_X32 U_g4176 ( .A(g2079), .ZN(g4176) );
INV_X32 U_g4179 ( .A(g2106), .ZN(g4179) );
INV_X32 U_g4182 ( .A(g2223), .ZN(g4182) );
INV_X32 U_g4185 ( .A(g2228), .ZN(g4185) );
INV_X32 U_g4188 ( .A(g2230), .ZN(g4188) );
INV_X32 U_g4191 ( .A(g2244), .ZN(g4191) );
INV_X32 U_g4194 ( .A(g2249), .ZN(g4194) );
INV_X32 U_g4197 ( .A(g2251), .ZN(g4197) );
INV_X32 U_I13366 ( .A(g2851), .ZN(I13366) );
INV_X32 U_g4200 ( .A(I13366), .ZN(g4200) );
INV_X32 U_g4201 ( .A(g2851), .ZN(g4201) );
INV_X32 U_g4202 ( .A(g42), .ZN(g4202) );
INV_X32 U_g4203 ( .A(g20), .ZN(g4203) );
INV_X32 U_g4204 ( .A(g3188), .ZN(g4204) );
INV_X32 U_g4205 ( .A(g131), .ZN(g4205) );
INV_X32 U_g4208 ( .A(g133), .ZN(g4208) );
INV_X32 U_g4211 ( .A(g159), .ZN(g4211) );
INV_X32 U_g4214 ( .A(g164), .ZN(g4214) );
INV_X32 U_g4217 ( .A(g354), .ZN(g4217) );
INV_X32 U_g4220 ( .A(g423), .ZN(g4220) );
INV_X32 U_g4221 ( .A(g426), .ZN(g4221) );
INV_X32 U_g4224 ( .A(g429), .ZN(g4224) );
INV_X32 U_g4225 ( .A(g701), .ZN(g4225) );
INV_X32 U_g4228 ( .A(g706), .ZN(g4228) );
INV_X32 U_g4231 ( .A(g708), .ZN(g4231) );
INV_X32 U_g4234 ( .A(g818), .ZN(g4234) );
INV_X32 U_g4237 ( .A(g844), .ZN(g4237) );
INV_X32 U_g4240 ( .A(g849), .ZN(g4240) );
INV_X32 U_g4243 ( .A(g851), .ZN(g4243) );
INV_X32 U_g4246 ( .A(g865), .ZN(g4246) );
INV_X32 U_g4249 ( .A(g1101), .ZN(g4249) );
INV_X32 U_g4250 ( .A(g1107), .ZN(g4250) );
INV_X32 U_g4251 ( .A(g1115), .ZN(g4251) );
INV_X32 U_g4254 ( .A(g1384), .ZN(g4254) );
INV_X32 U_g4257 ( .A(g1389), .ZN(g4257) );
INV_X32 U_g4260 ( .A(g1391), .ZN(g4260) );
INV_X32 U_g4263 ( .A(g1411), .ZN(g4263) );
INV_X32 U_g4266 ( .A(g1535), .ZN(g4266) );
INV_X32 U_g4269 ( .A(g1540), .ZN(g4269) );
INV_X32 U_g4272 ( .A(g1542), .ZN(g4272) );
INV_X32 U_g4275 ( .A(g1556), .ZN(g4275) );
INV_X32 U_g4278 ( .A(g1561), .ZN(g4278) );
INV_X32 U_g4281 ( .A(g1792), .ZN(g4281) );
INV_X32 U_g4282 ( .A(g1798), .ZN(g4282) );
INV_X32 U_g4283 ( .A(g1808), .ZN(g4283) );
INV_X32 U_g4286 ( .A(g2080), .ZN(g4286) );
INV_X32 U_g4289 ( .A(g2082), .ZN(g4289) );
INV_X32 U_g4292 ( .A(g2107), .ZN(g4292) );
INV_X32 U_g4295 ( .A(g2226), .ZN(g4295) );
INV_X32 U_g4298 ( .A(g2231), .ZN(g4298) );
INV_X32 U_g4301 ( .A(g2233), .ZN(g4301) );
INV_X32 U_g4304 ( .A(g2247), .ZN(g4304) );
INV_X32 U_g4307 ( .A(g2252), .ZN(g4307) );
INV_X32 U_g4310 ( .A(g2254), .ZN(g4310) );
INV_X32 U_g4313 ( .A(g2483), .ZN(g4313) );
INV_X32 U_g4314 ( .A(g2530), .ZN(g4314) );
INV_X32 U_g4315 ( .A(g2773), .ZN(g4315) );
INV_X32 U_g4318 ( .A(g2800), .ZN(g4318) );
INV_X32 U_I13417 ( .A(g2839), .ZN(I13417) );
INV_X32 U_g4321 ( .A(I13417), .ZN(g4321) );
INV_X32 U_g4322 ( .A(g2839), .ZN(g4322) );
INV_X32 U_I13421 ( .A(g2867), .ZN(I13421) );
INV_X32 U_g4323 ( .A(I13421), .ZN(g4323) );
INV_X32 U_g4324 ( .A(g2867), .ZN(g4324) );
INV_X32 U_g4325 ( .A(g36), .ZN(g4325) );
INV_X32 U_g4326 ( .A(g181), .ZN(g4326) );
INV_X32 U_g4329 ( .A(g129), .ZN(g4329) );
INV_X32 U_g4332 ( .A(g134), .ZN(g4332) );
INV_X32 U_g4335 ( .A(g162), .ZN(g4335) );
INV_X32 U_I13430 ( .A(g101), .ZN(I13430) );
INV_X32 U_g4338 ( .A(I13430), .ZN(g4338) );
INV_X32 U_I13433 ( .A(g105), .ZN(I13433) );
INV_X32 U_g4339 ( .A(I13433), .ZN(g4339) );
INV_X32 U_g4340 ( .A(g343), .ZN(g4340) );
INV_X32 U_g4343 ( .A(g369), .ZN(g4343) );
INV_X32 U_g4346 ( .A(g432), .ZN(g4346) );
INV_X32 U_g4347 ( .A(g438), .ZN(g4347) );
INV_X32 U_g4348 ( .A(g704), .ZN(g4348) );
INV_X32 U_g4351 ( .A(g709), .ZN(g4351) );
INV_X32 U_g4354 ( .A(g711), .ZN(g4354) );
INV_X32 U_g4357 ( .A(g729), .ZN(g4357) );
INV_X32 U_g4360 ( .A(g819), .ZN(g4360) );
INV_X32 U_g4363 ( .A(g821), .ZN(g4363) );
INV_X32 U_g4366 ( .A(g847), .ZN(g4366) );
INV_X32 U_g4369 ( .A(g852), .ZN(g4369) );
INV_X32 U_g4372 ( .A(g1041), .ZN(g4372) );
INV_X32 U_g4375 ( .A(g1110), .ZN(g4375) );
INV_X32 U_g4376 ( .A(g1113), .ZN(g4376) );
INV_X32 U_g4379 ( .A(g1116), .ZN(g4379) );
INV_X32 U_g4380 ( .A(g1387), .ZN(g4380) );
INV_X32 U_g4383 ( .A(g1392), .ZN(g4383) );
INV_X32 U_g4386 ( .A(g1394), .ZN(g4386) );
INV_X32 U_g4389 ( .A(g1512), .ZN(g4389) );
INV_X32 U_g4392 ( .A(g1538), .ZN(g4392) );
INV_X32 U_g4395 ( .A(g1543), .ZN(g4395) );
INV_X32 U_g4398 ( .A(g1545), .ZN(g4398) );
INV_X32 U_g4401 ( .A(g1559), .ZN(g4401) );
INV_X32 U_g4404 ( .A(g1795), .ZN(g4404) );
INV_X32 U_g4405 ( .A(g1801), .ZN(g4405) );
INV_X32 U_g4406 ( .A(g1809), .ZN(g4406) );
INV_X32 U_g4409 ( .A(g2078), .ZN(g4409) );
INV_X32 U_g4412 ( .A(g2083), .ZN(g4412) );
INV_X32 U_g4415 ( .A(g2085), .ZN(g4415) );
INV_X32 U_g4418 ( .A(g2105), .ZN(g4418) );
INV_X32 U_g4421 ( .A(g2229), .ZN(g4421) );
INV_X32 U_g4424 ( .A(g2234), .ZN(g4424) );
INV_X32 U_g4427 ( .A(g2236), .ZN(g4427) );
INV_X32 U_g4430 ( .A(g2250), .ZN(g4430) );
INV_X32 U_g4433 ( .A(g2255), .ZN(g4433) );
INV_X32 U_g4436 ( .A(g2486), .ZN(g4436) );
INV_X32 U_g4437 ( .A(g2492), .ZN(g4437) );
INV_X32 U_g4438 ( .A(g2502), .ZN(g4438) );
INV_X32 U_g4441 ( .A(g2774), .ZN(g4441) );
INV_X32 U_g4444 ( .A(g2776), .ZN(g4444) );
INV_X32 U_g4447 ( .A(g2801), .ZN(g4447) );
INV_X32 U_I13478 ( .A(g2854), .ZN(I13478) );
INV_X32 U_g4450 ( .A(I13478), .ZN(g4450) );
INV_X32 U_g4451 ( .A(g2854), .ZN(g4451) );
INV_X32 U_g4452 ( .A(g17), .ZN(g4452) );
INV_X32 U_g4453 ( .A(g132), .ZN(g4453) );
INV_X32 U_g4456 ( .A(g309), .ZN(g4456) );
INV_X32 U_g4465 ( .A(g346), .ZN(g4465) );
INV_X32 U_g4468 ( .A(g358), .ZN(g4468) );
INV_X32 U_g4471 ( .A(g384), .ZN(g4471) );
INV_X32 U_g4474 ( .A(g435), .ZN(g4474) );
INV_X32 U_g4475 ( .A(g441), .ZN(g4475) );
INV_X32 U_g4476 ( .A(g576), .ZN(g4476) );
INV_X32 U_g4479 ( .A(g587), .ZN(g4479) );
INV_X32 U_g4480 ( .A(g707), .ZN(g4480) );
INV_X32 U_g4483 ( .A(g712), .ZN(g4483) );
INV_X32 U_g4486 ( .A(g714), .ZN(g4486) );
INV_X32 U_g4489 ( .A(g730), .ZN(g4489) );
INV_X32 U_g4492 ( .A(g732), .ZN(g4492) );
INV_X32 U_g4495 ( .A(g869), .ZN(g4495) );
INV_X32 U_g4498 ( .A(g817), .ZN(g4498) );
INV_X32 U_g4501 ( .A(g822), .ZN(g4501) );
INV_X32 U_g4504 ( .A(g850), .ZN(g4504) );
INV_X32 U_I13501 ( .A(g789), .ZN(I13501) );
INV_X32 U_g4507 ( .A(I13501), .ZN(g4507) );
INV_X32 U_I13504 ( .A(g793), .ZN(I13504) );
INV_X32 U_g4508 ( .A(I13504), .ZN(g4508) );
INV_X32 U_g4509 ( .A(g1030), .ZN(g4509) );
INV_X32 U_g4512 ( .A(g1056), .ZN(g4512) );
INV_X32 U_g4515 ( .A(g1119), .ZN(g4515) );
INV_X32 U_g4516 ( .A(g1125), .ZN(g4516) );
INV_X32 U_g4517 ( .A(g1390), .ZN(g4517) );
INV_X32 U_g4520 ( .A(g1395), .ZN(g4520) );
INV_X32 U_g4523 ( .A(g1397), .ZN(g4523) );
INV_X32 U_g4526 ( .A(g1415), .ZN(g4526) );
INV_X32 U_g4529 ( .A(g1513), .ZN(g4529) );
INV_X32 U_g4532 ( .A(g1515), .ZN(g4532) );
INV_X32 U_g4535 ( .A(g1541), .ZN(g4535) );
INV_X32 U_g4538 ( .A(g1546), .ZN(g4538) );
INV_X32 U_g4541 ( .A(g1735), .ZN(g4541) );
INV_X32 U_g4544 ( .A(g1804), .ZN(g4544) );
INV_X32 U_g4545 ( .A(g1807), .ZN(g4545) );
INV_X32 U_g4548 ( .A(g1810), .ZN(g4548) );
INV_X32 U_g4549 ( .A(g2081), .ZN(g4549) );
INV_X32 U_g4552 ( .A(g2086), .ZN(g4552) );
INV_X32 U_g4555 ( .A(g2088), .ZN(g4555) );
INV_X32 U_g4558 ( .A(g2206), .ZN(g4558) );
INV_X32 U_g4561 ( .A(g2232), .ZN(g4561) );
INV_X32 U_g4564 ( .A(g2237), .ZN(g4564) );
INV_X32 U_g4567 ( .A(g2239), .ZN(g4567) );
INV_X32 U_g4570 ( .A(g2253), .ZN(g4570) );
INV_X32 U_g4573 ( .A(g2489), .ZN(g4573) );
INV_X32 U_g4574 ( .A(g2495), .ZN(g4574) );
INV_X32 U_g4575 ( .A(g2503), .ZN(g4575) );
INV_X32 U_g4578 ( .A(g2772), .ZN(g4578) );
INV_X32 U_g4581 ( .A(g2777), .ZN(g4581) );
INV_X32 U_g4584 ( .A(g2779), .ZN(g4584) );
INV_X32 U_g4587 ( .A(g2799), .ZN(g4587) );
INV_X32 U_I13538 ( .A(g2870), .ZN(I13538) );
INV_X32 U_g4590 ( .A(I13538), .ZN(g4590) );
INV_X32 U_g4591 ( .A(g2870), .ZN(g4591) );
INV_X32 U_g4592 ( .A(g361), .ZN(g4592) );
INV_X32 U_g4595 ( .A(g373), .ZN(g4595) );
INV_X32 U_g4598 ( .A(g398), .ZN(g4598) );
INV_X32 U_g4601 ( .A(g444), .ZN(g4601) );
INV_X32 U_g4602 ( .A(g525), .ZN(g4602) );
INV_X32 U_g4603 ( .A(g577), .ZN(g4603) );
INV_X32 U_g4606 ( .A(g579), .ZN(g4606) );
INV_X32 U_g4609 ( .A(g590), .ZN(g4609) );
INV_X32 U_g4610 ( .A(g596), .ZN(g4610) );
INV_X32 U_g4611 ( .A(g710), .ZN(g4611) );
INV_X32 U_g4614 ( .A(g715), .ZN(g4614) );
INV_X32 U_g4617 ( .A(g717), .ZN(g4617) );
INV_X32 U_g4620 ( .A(g728), .ZN(g4620) );
INV_X32 U_g4623 ( .A(g733), .ZN(g4623) );
INV_X32 U_g4626 ( .A(g735), .ZN(g4626) );
INV_X32 U_g4629 ( .A(g820), .ZN(g4629) );
INV_X32 U_g4632 ( .A(g996), .ZN(g4632) );
INV_X32 U_g4641 ( .A(g1033), .ZN(g4641) );
INV_X32 U_g4644 ( .A(g1045), .ZN(g4644) );
INV_X32 U_g4647 ( .A(g1071), .ZN(g4647) );
INV_X32 U_g4650 ( .A(g1122), .ZN(g4650) );
INV_X32 U_g4651 ( .A(g1128), .ZN(g4651) );
INV_X32 U_g4652 ( .A(g1262), .ZN(g4652) );
INV_X32 U_g4655 ( .A(g1273), .ZN(g4655) );
INV_X32 U_g4656 ( .A(g1393), .ZN(g4656) );
INV_X32 U_g4659 ( .A(g1398), .ZN(g4659) );
INV_X32 U_g4662 ( .A(g1400), .ZN(g4662) );
INV_X32 U_g4665 ( .A(g1416), .ZN(g4665) );
INV_X32 U_g4668 ( .A(g1418), .ZN(g4668) );
INV_X32 U_g4671 ( .A(g1563), .ZN(g4671) );
INV_X32 U_g4674 ( .A(g1511), .ZN(g4674) );
INV_X32 U_g4677 ( .A(g1516), .ZN(g4677) );
INV_X32 U_g4680 ( .A(g1544), .ZN(g4680) );
INV_X32 U_I13575 ( .A(g1476), .ZN(I13575) );
INV_X32 U_g4683 ( .A(I13575), .ZN(g4683) );
INV_X32 U_I13578 ( .A(g1481), .ZN(I13578) );
INV_X32 U_g4684 ( .A(I13578), .ZN(g4684) );
INV_X32 U_g4685 ( .A(g1724), .ZN(g4685) );
INV_X32 U_g4688 ( .A(g1750), .ZN(g4688) );
INV_X32 U_g4691 ( .A(g1813), .ZN(g4691) );
INV_X32 U_g4692 ( .A(g1819), .ZN(g4692) );
INV_X32 U_g4693 ( .A(g2084), .ZN(g4693) );
INV_X32 U_g4696 ( .A(g2089), .ZN(g4696) );
INV_X32 U_g4699 ( .A(g2091), .ZN(g4699) );
INV_X32 U_g4702 ( .A(g2109), .ZN(g4702) );
INV_X32 U_g4705 ( .A(g2207), .ZN(g4705) );
INV_X32 U_g4708 ( .A(g2209), .ZN(g4708) );
INV_X32 U_g4711 ( .A(g2235), .ZN(g4711) );
INV_X32 U_g4714 ( .A(g2240), .ZN(g4714) );
INV_X32 U_g4717 ( .A(g2429), .ZN(g4717) );
INV_X32 U_g4720 ( .A(g2498), .ZN(g4720) );
INV_X32 U_g4721 ( .A(g2501), .ZN(g4721) );
INV_X32 U_g4724 ( .A(g2504), .ZN(g4724) );
INV_X32 U_g4725 ( .A(g2775), .ZN(g4725) );
INV_X32 U_g4728 ( .A(g2780), .ZN(g4728) );
INV_X32 U_g4731 ( .A(g2782), .ZN(g4731) );
INV_X32 U_g4734 ( .A(g11), .ZN(g4734) );
INV_X32 U_I13601 ( .A(g121), .ZN(I13601) );
INV_X32 U_g4735 ( .A(I13601), .ZN(g4735) );
INV_X32 U_I13604 ( .A(g125), .ZN(I13604) );
INV_X32 U_g4736 ( .A(I13604), .ZN(g4736) );
INV_X32 U_g4737 ( .A(g376), .ZN(g4737) );
INV_X32 U_g4740 ( .A(g388), .ZN(g4740) );
INV_X32 U_g4743 ( .A(g575), .ZN(g4743) );
INV_X32 U_g4746 ( .A(g580), .ZN(g4746) );
INV_X32 U_g4749 ( .A(g582), .ZN(g4749) );
INV_X32 U_g4752 ( .A(g593), .ZN(g4752) );
INV_X32 U_g4753 ( .A(g599), .ZN(g4753) );
INV_X32 U_g4754 ( .A(g713), .ZN(g4754) );
INV_X32 U_g4757 ( .A(g718), .ZN(g4757) );
INV_X32 U_g4760 ( .A(g720), .ZN(g4760) );
INV_X32 U_g4763 ( .A(g731), .ZN(g4763) );
INV_X32 U_g4766 ( .A(g736), .ZN(g4766) );
INV_X32 U_g4769 ( .A(g1048), .ZN(g4769) );
INV_X32 U_g4772 ( .A(g1060), .ZN(g4772) );
INV_X32 U_g4775 ( .A(g1085), .ZN(g4775) );
INV_X32 U_g4778 ( .A(g1131), .ZN(g4778) );
INV_X32 U_g4779 ( .A(g1211), .ZN(g4779) );
INV_X32 U_g4780 ( .A(g1263), .ZN(g4780) );
INV_X32 U_g4783 ( .A(g1265), .ZN(g4783) );
INV_X32 U_g4786 ( .A(g1276), .ZN(g4786) );
INV_X32 U_g4787 ( .A(g1282), .ZN(g4787) );
INV_X32 U_g4788 ( .A(g1396), .ZN(g4788) );
INV_X32 U_g4791 ( .A(g1401), .ZN(g4791) );
INV_X32 U_g4794 ( .A(g1403), .ZN(g4794) );
INV_X32 U_g4797 ( .A(g1414), .ZN(g4797) );
INV_X32 U_g4800 ( .A(g1419), .ZN(g4800) );
INV_X32 U_g4803 ( .A(g1421), .ZN(g4803) );
INV_X32 U_g4806 ( .A(g1514), .ZN(g4806) );
INV_X32 U_g4809 ( .A(g1690), .ZN(g4809) );
INV_X32 U_g4818 ( .A(g1727), .ZN(g4818) );
INV_X32 U_g4821 ( .A(g1739), .ZN(g4821) );
INV_X32 U_g4824 ( .A(g1765), .ZN(g4824) );
INV_X32 U_g4827 ( .A(g1816), .ZN(g4827) );
INV_X32 U_g4828 ( .A(g1822), .ZN(g4828) );
INV_X32 U_g4829 ( .A(g1956), .ZN(g4829) );
INV_X32 U_g4832 ( .A(g1967), .ZN(g4832) );
INV_X32 U_g4833 ( .A(g2087), .ZN(g4833) );
INV_X32 U_g4836 ( .A(g2092), .ZN(g4836) );
INV_X32 U_g4839 ( .A(g2094), .ZN(g4839) );
INV_X32 U_g4842 ( .A(g2110), .ZN(g4842) );
INV_X32 U_g4845 ( .A(g2112), .ZN(g4845) );
INV_X32 U_g4848 ( .A(g2257), .ZN(g4848) );
INV_X32 U_g4851 ( .A(g2205), .ZN(g4851) );
INV_X32 U_g4854 ( .A(g2210), .ZN(g4854) );
INV_X32 U_g4857 ( .A(g2238), .ZN(g4857) );
INV_X32 U_I13652 ( .A(g2170), .ZN(I13652) );
INV_X32 U_g4860 ( .A(I13652), .ZN(g4860) );
INV_X32 U_I13655 ( .A(g2175), .ZN(I13655) );
INV_X32 U_g4861 ( .A(I13655), .ZN(g4861) );
INV_X32 U_g4862 ( .A(g2418), .ZN(g4862) );
INV_X32 U_g4865 ( .A(g2444), .ZN(g4865) );
INV_X32 U_g4868 ( .A(g2507), .ZN(g4868) );
INV_X32 U_g4869 ( .A(g2513), .ZN(g4869) );
INV_X32 U_g4870 ( .A(g2778), .ZN(g4870) );
INV_X32 U_g4873 ( .A(g2783), .ZN(g4873) );
INV_X32 U_g4876 ( .A(g2785), .ZN(g4876) );
INV_X32 U_g4879 ( .A(g2803), .ZN(g4879) );
INV_X32 U_g4882 ( .A(g391), .ZN(g4882) );
INV_X32 U_g4885 ( .A(g448), .ZN(g4885) );
INV_X32 U_g4888 ( .A(g578), .ZN(g4888) );
INV_X32 U_g4891 ( .A(g583), .ZN(g4891) );
INV_X32 U_g4894 ( .A(g585), .ZN(g4894) );
INV_X32 U_g4897 ( .A(g602), .ZN(g4897) );
INV_X32 U_g4898 ( .A(g605), .ZN(g4898) );
INV_X32 U_g4899 ( .A(g716), .ZN(g4899) );
INV_X32 U_g4902 ( .A(g721), .ZN(g4902) );
INV_X32 U_g4905 ( .A(g723), .ZN(g4905) );
INV_X32 U_g4908 ( .A(g734), .ZN(g4908) );
INV_X32 U_I13677 ( .A(g809), .ZN(I13677) );
INV_X32 U_g4911 ( .A(I13677), .ZN(g4911) );
INV_X32 U_I13680 ( .A(g813), .ZN(I13680) );
INV_X32 U_g4912 ( .A(I13680), .ZN(g4912) );
INV_X32 U_g4913 ( .A(g1063), .ZN(g4913) );
INV_X32 U_g4916 ( .A(g1075), .ZN(g4916) );
INV_X32 U_g4919 ( .A(g1261), .ZN(g4919) );
INV_X32 U_g4922 ( .A(g1266), .ZN(g4922) );
INV_X32 U_g4925 ( .A(g1268), .ZN(g4925) );
INV_X32 U_g4928 ( .A(g1279), .ZN(g4928) );
INV_X32 U_g4929 ( .A(g1285), .ZN(g4929) );
INV_X32 U_g4930 ( .A(g1399), .ZN(g4930) );
INV_X32 U_g4933 ( .A(g1404), .ZN(g4933) );
INV_X32 U_g4936 ( .A(g1406), .ZN(g4936) );
INV_X32 U_g4939 ( .A(g1417), .ZN(g4939) );
INV_X32 U_g4942 ( .A(g1422), .ZN(g4942) );
INV_X32 U_g4945 ( .A(g1742), .ZN(g4945) );
INV_X32 U_g4948 ( .A(g1754), .ZN(g4948) );
INV_X32 U_g4951 ( .A(g1779), .ZN(g4951) );
INV_X32 U_g4954 ( .A(g1825), .ZN(g4954) );
INV_X32 U_g4955 ( .A(g1905), .ZN(g4955) );
INV_X32 U_g4956 ( .A(g1957), .ZN(g4956) );
INV_X32 U_g4959 ( .A(g1959), .ZN(g4959) );
INV_X32 U_g4962 ( .A(g1970), .ZN(g4962) );
INV_X32 U_g4963 ( .A(g1976), .ZN(g4963) );
INV_X32 U_g4964 ( .A(g2090), .ZN(g4964) );
INV_X32 U_g4967 ( .A(g2095), .ZN(g4967) );
INV_X32 U_g4970 ( .A(g2097), .ZN(g4970) );
INV_X32 U_g4973 ( .A(g2108), .ZN(g4973) );
INV_X32 U_g4976 ( .A(g2113), .ZN(g4976) );
INV_X32 U_g4979 ( .A(g2115), .ZN(g4979) );
INV_X32 U_g4982 ( .A(g2208), .ZN(g4982) );
INV_X32 U_g4985 ( .A(g2384), .ZN(g4985) );
INV_X32 U_g4994 ( .A(g2421), .ZN(g4994) );
INV_X32 U_g4997 ( .A(g2433), .ZN(g4997) );
INV_X32 U_g5000 ( .A(g2459), .ZN(g5000) );
INV_X32 U_g5003 ( .A(g2510), .ZN(g5003) );
INV_X32 U_g5004 ( .A(g2516), .ZN(g5004) );
INV_X32 U_g5005 ( .A(g2650), .ZN(g5005) );
INV_X32 U_g5008 ( .A(g2661), .ZN(g5008) );
INV_X32 U_g5009 ( .A(g2781), .ZN(g5009) );
INV_X32 U_g5012 ( .A(g2786), .ZN(g5012) );
INV_X32 U_g5015 ( .A(g2788), .ZN(g5015) );
INV_X32 U_g5018 ( .A(g2804), .ZN(g5018) );
INV_X32 U_g5021 ( .A(g2806), .ZN(g5021) );
INV_X32 U_g5024 ( .A(g449), .ZN(g5024) );
INV_X32 U_g5027 ( .A(g581), .ZN(g5027) );
INV_X32 U_g5030 ( .A(g586), .ZN(g5030) );
INV_X32 U_g5033 ( .A(g608), .ZN(g5033) );
INV_X32 U_g5034 ( .A(g614), .ZN(g5034) );
INV_X32 U_g5035 ( .A(g719), .ZN(g5035) );
INV_X32 U_g5038 ( .A(g724), .ZN(g5038) );
INV_X32 U_g5041 ( .A(g1078), .ZN(g5041) );
INV_X32 U_g5044 ( .A(g1135), .ZN(g5044) );
INV_X32 U_g5047 ( .A(g1264), .ZN(g5047) );
INV_X32 U_g5050 ( .A(g1269), .ZN(g5050) );
INV_X32 U_g5053 ( .A(g1271), .ZN(g5053) );
INV_X32 U_g5056 ( .A(g1288), .ZN(g5056) );
INV_X32 U_g5057 ( .A(g1291), .ZN(g5057) );
INV_X32 U_g5058 ( .A(g1402), .ZN(g5058) );
INV_X32 U_g5061 ( .A(g1407), .ZN(g5061) );
INV_X32 U_g5064 ( .A(g1409), .ZN(g5064) );
INV_X32 U_g5067 ( .A(g1420), .ZN(g5067) );
INV_X32 U_I13742 ( .A(g1501), .ZN(I13742) );
INV_X32 U_g5070 ( .A(I13742), .ZN(g5070) );
INV_X32 U_I13745 ( .A(g1506), .ZN(I13745) );
INV_X32 U_g5071 ( .A(I13745), .ZN(g5071) );
INV_X32 U_g5072 ( .A(g1757), .ZN(g5072) );
INV_X32 U_g5075 ( .A(g1769), .ZN(g5075) );
INV_X32 U_g5078 ( .A(g1955), .ZN(g5078) );
INV_X32 U_g5081 ( .A(g1960), .ZN(g5081) );
INV_X32 U_g5084 ( .A(g1962), .ZN(g5084) );
INV_X32 U_g5087 ( .A(g1973), .ZN(g5087) );
INV_X32 U_g5088 ( .A(g1979), .ZN(g5088) );
INV_X32 U_g5089 ( .A(g2093), .ZN(g5089) );
INV_X32 U_g5092 ( .A(g2098), .ZN(g5092) );
INV_X32 U_g5095 ( .A(g2100), .ZN(g5095) );
INV_X32 U_g5098 ( .A(g2111), .ZN(g5098) );
INV_X32 U_g5101 ( .A(g2116), .ZN(g5101) );
INV_X32 U_g5104 ( .A(g2436), .ZN(g5104) );
INV_X32 U_g5107 ( .A(g2448), .ZN(g5107) );
INV_X32 U_g5110 ( .A(g2473), .ZN(g5110) );
INV_X32 U_g5113 ( .A(g2519), .ZN(g5113) );
INV_X32 U_g5114 ( .A(g2599), .ZN(g5114) );
INV_X32 U_g5115 ( .A(g2651), .ZN(g5115) );
INV_X32 U_g5118 ( .A(g2653), .ZN(g5118) );
INV_X32 U_g5121 ( .A(g2664), .ZN(g5121) );
INV_X32 U_g5122 ( .A(g2670), .ZN(g5122) );
INV_X32 U_g5123 ( .A(g2784), .ZN(g5123) );
INV_X32 U_g5126 ( .A(g2789), .ZN(g5126) );
INV_X32 U_g5129 ( .A(g2791), .ZN(g5129) );
INV_X32 U_g5132 ( .A(g2802), .ZN(g5132) );
INV_X32 U_g5135 ( .A(g2807), .ZN(g5135) );
INV_X32 U_g5138 ( .A(g2809), .ZN(g5138) );
INV_X32 U_I13775 ( .A(g109), .ZN(I13775) );
INV_X32 U_g5141 ( .A(I13775), .ZN(g5141) );
INV_X32 U_g5142 ( .A(g447), .ZN(g5142) );
INV_X32 U_g5145 ( .A(g584), .ZN(g5145) );
INV_X32 U_g5148 ( .A(g611), .ZN(g5148) );
INV_X32 U_g5149 ( .A(g617), .ZN(g5149) );
INV_X32 U_g5150 ( .A(g722), .ZN(g5150) );
INV_X32 U_g5153 ( .A(g1136), .ZN(g5153) );
INV_X32 U_g5156 ( .A(g1267), .ZN(g5156) );
INV_X32 U_g5159 ( .A(g1272), .ZN(g5159) );
INV_X32 U_g5162 ( .A(g1294), .ZN(g5162) );
INV_X32 U_g5163 ( .A(g1300), .ZN(g5163) );
INV_X32 U_g5164 ( .A(g1405), .ZN(g5164) );
INV_X32 U_g5167 ( .A(g1410), .ZN(g5167) );
INV_X32 U_g5170 ( .A(g1772), .ZN(g5170) );
INV_X32 U_g5173 ( .A(g1829), .ZN(g5173) );
INV_X32 U_g5176 ( .A(g1958), .ZN(g5176) );
INV_X32 U_g5179 ( .A(g1963), .ZN(g5179) );
INV_X32 U_g5182 ( .A(g1965), .ZN(g5182) );
INV_X32 U_g5185 ( .A(g1982), .ZN(g5185) );
INV_X32 U_g5186 ( .A(g1985), .ZN(g5186) );
INV_X32 U_g5187 ( .A(g2096), .ZN(g5187) );
INV_X32 U_g5190 ( .A(g2101), .ZN(g5190) );
INV_X32 U_g5193 ( .A(g2103), .ZN(g5193) );
INV_X32 U_g5196 ( .A(g2114), .ZN(g5196) );
INV_X32 U_I13801 ( .A(g2195), .ZN(I13801) );
INV_X32 U_g5199 ( .A(I13801), .ZN(g5199) );
INV_X32 U_I13804 ( .A(g2200), .ZN(I13804) );
INV_X32 U_g5200 ( .A(I13804), .ZN(g5200) );
INV_X32 U_g5201 ( .A(g2451), .ZN(g5201) );
INV_X32 U_g5204 ( .A(g2463), .ZN(g5204) );
INV_X32 U_g5207 ( .A(g2649), .ZN(g5207) );
INV_X32 U_g5210 ( .A(g2654), .ZN(g5210) );
INV_X32 U_g5213 ( .A(g2656), .ZN(g5213) );
INV_X32 U_g5216 ( .A(g2667), .ZN(g5216) );
INV_X32 U_g5217 ( .A(g2673), .ZN(g5217) );
INV_X32 U_g5218 ( .A(g2787), .ZN(g5218) );
INV_X32 U_g5221 ( .A(g2792), .ZN(g5221) );
INV_X32 U_g5224 ( .A(g2794), .ZN(g5224) );
INV_X32 U_g5227 ( .A(g2805), .ZN(g5227) );
INV_X32 U_g5230 ( .A(g2810), .ZN(g5230) );
INV_X32 U_g5233 ( .A(g620), .ZN(g5233) );
INV_X32 U_I13820 ( .A(g797), .ZN(I13820) );
INV_X32 U_g5234 ( .A(I13820), .ZN(g5234) );
INV_X32 U_g5235 ( .A(g1134), .ZN(g5235) );
INV_X32 U_g5238 ( .A(g1270), .ZN(g5238) );
INV_X32 U_g5241 ( .A(g1297), .ZN(g5241) );
INV_X32 U_g5242 ( .A(g1303), .ZN(g5242) );
INV_X32 U_g5243 ( .A(g1408), .ZN(g5243) );
INV_X32 U_g5246 ( .A(g1830), .ZN(g5246) );
INV_X32 U_g5249 ( .A(g1961), .ZN(g5249) );
INV_X32 U_g5252 ( .A(g1966), .ZN(g5252) );
INV_X32 U_g5255 ( .A(g1988), .ZN(g5255) );
INV_X32 U_g5256 ( .A(g1994), .ZN(g5256) );
INV_X32 U_g5257 ( .A(g2099), .ZN(g5257) );
INV_X32 U_g5260 ( .A(g2104), .ZN(g5260) );
INV_X32 U_g5263 ( .A(g2466), .ZN(g5263) );
INV_X32 U_g5266 ( .A(g2523), .ZN(g5266) );
INV_X32 U_g5269 ( .A(g2652), .ZN(g5269) );
INV_X32 U_g5272 ( .A(g2657), .ZN(g5272) );
INV_X32 U_g5275 ( .A(g2659), .ZN(g5275) );
INV_X32 U_g5278 ( .A(g2676), .ZN(g5278) );
INV_X32 U_g5279 ( .A(g2679), .ZN(g5279) );
INV_X32 U_g5280 ( .A(g2790), .ZN(g5280) );
INV_X32 U_g5283 ( .A(g2795), .ZN(g5283) );
INV_X32 U_g5286 ( .A(g2797), .ZN(g5286) );
INV_X32 U_g5289 ( .A(g2808), .ZN(g5289) );
INV_X32 U_g5292 ( .A(g2857), .ZN(g5292) );
INV_X32 U_g5293 ( .A(g738), .ZN(g5293) );
INV_X32 U_g5296 ( .A(g1306), .ZN(g5296) );
INV_X32 U_I13849 ( .A(g1486), .ZN(I13849) );
INV_X32 U_g5297 ( .A(I13849), .ZN(g5297) );
INV_X32 U_g5298 ( .A(g1828), .ZN(g5298) );
INV_X32 U_g5301 ( .A(g1964), .ZN(g5301) );
INV_X32 U_g5304 ( .A(g1991), .ZN(g5304) );
INV_X32 U_g5305 ( .A(g1997), .ZN(g5305) );
INV_X32 U_g5306 ( .A(g2102), .ZN(g5306) );
INV_X32 U_g5309 ( .A(g2524), .ZN(g5309) );
INV_X32 U_g5312 ( .A(g2655), .ZN(g5312) );
INV_X32 U_g5315 ( .A(g2660), .ZN(g5315) );
INV_X32 U_g5318 ( .A(g2682), .ZN(g5318) );
INV_X32 U_g5319 ( .A(g2688), .ZN(g5319) );
INV_X32 U_g5320 ( .A(g2793), .ZN(g5320) );
INV_X32 U_g5323 ( .A(g2798), .ZN(g5323) );
INV_X32 U_g5326 ( .A(g2873), .ZN(g5326) );
INV_X32 U_g5327 ( .A(g739), .ZN(g5327) );
INV_X32 U_g5330 ( .A(g1424), .ZN(g5330) );
INV_X32 U_g5333 ( .A(g2000), .ZN(g5333) );
INV_X32 U_I13868 ( .A(g2180), .ZN(I13868) );
INV_X32 U_g5334 ( .A(I13868), .ZN(g5334) );
INV_X32 U_g5335 ( .A(g2522), .ZN(g5335) );
INV_X32 U_g5338 ( .A(g2658), .ZN(g5338) );
INV_X32 U_g5341 ( .A(g2685), .ZN(g5341) );
INV_X32 U_g5342 ( .A(g2691), .ZN(g5342) );
INV_X32 U_g5343 ( .A(g2796), .ZN(g5343) );
INV_X32 U_g5346 ( .A(g3106), .ZN(g5346) );
INV_X32 U_g5349 ( .A(g2877), .ZN(g5349) );
INV_X32 U_g5352 ( .A(g737), .ZN(g5352) );
INV_X32 U_g5355 ( .A(g1425), .ZN(g5355) );
INV_X32 U_g5358 ( .A(g2118), .ZN(g5358) );
INV_X32 U_g5361 ( .A(g2694), .ZN(g5361) );
INV_X32 U_g5362 ( .A(g2817), .ZN(g5362) );
INV_X32 U_g5363 ( .A(g3107), .ZN(g5363) );
INV_X32 U_g5366 ( .A(g2878), .ZN(g5366) );
INV_X32 U_g5369 ( .A(g1423), .ZN(g5369) );
INV_X32 U_g5372 ( .A(g2119), .ZN(g5372) );
INV_X32 U_g5375 ( .A(g2812), .ZN(g5375) );
INV_X32 U_g5378 ( .A(g2933), .ZN(g5378) );
INV_X32 U_g5379 ( .A(g3108), .ZN(g5379) );
INV_X32 U_g5382 ( .A(g2117), .ZN(g5382) );
INV_X32 U_g5385 ( .A(g2813), .ZN(g5385) );
INV_X32 U_I13892 ( .A(g3040), .ZN(I13892) );
INV_X32 U_g5388 ( .A(I13892), .ZN(g5388) );
INV_X32 U_g5389 ( .A(g3040), .ZN(g5389) );
INV_X32 U_I13896 ( .A(g343), .ZN(I13896) );
INV_X32 U_g5390 ( .A(I13896), .ZN(g5390) );
INV_X32 U_g5391 ( .A(g2811), .ZN(g5391) );
INV_X32 U_g5394 ( .A(g3054), .ZN(g5394) );
INV_X32 U_I13901 ( .A(g346), .ZN(I13901) );
INV_X32 U_g5395 ( .A(I13901), .ZN(g5395) );
INV_X32 U_I13904 ( .A(g358), .ZN(I13904) );
INV_X32 U_g5396 ( .A(I13904), .ZN(g5396) );
INV_X32 U_I13907 ( .A(g1030), .ZN(I13907) );
INV_X32 U_g5397 ( .A(I13907), .ZN(g5397) );
INV_X32 U_I13910 ( .A(g361), .ZN(I13910) );
INV_X32 U_g5398 ( .A(I13910), .ZN(g5398) );
INV_X32 U_I13913 ( .A(g373), .ZN(I13913) );
INV_X32 U_g5399 ( .A(I13913), .ZN(g5399) );
INV_X32 U_I13916 ( .A(g1033), .ZN(I13916) );
INV_X32 U_g5400 ( .A(I13916), .ZN(g5400) );
INV_X32 U_I13919 ( .A(g1045), .ZN(I13919) );
INV_X32 U_g5401 ( .A(I13919), .ZN(g5401) );
INV_X32 U_I13922 ( .A(g1724), .ZN(I13922) );
INV_X32 U_g5402 ( .A(I13922), .ZN(g5402) );
INV_X32 U_I13925 ( .A(g376), .ZN(I13925) );
INV_X32 U_g5403 ( .A(I13925), .ZN(g5403) );
INV_X32 U_I13928 ( .A(g388), .ZN(I13928) );
INV_X32 U_g5404 ( .A(I13928), .ZN(g5404) );
INV_X32 U_I13931 ( .A(g1048), .ZN(I13931) );
INV_X32 U_g5405 ( .A(I13931), .ZN(g5405) );
INV_X32 U_I13934 ( .A(g1060), .ZN(I13934) );
INV_X32 U_g5406 ( .A(I13934), .ZN(g5406) );
INV_X32 U_I13937 ( .A(g1727), .ZN(I13937) );
INV_X32 U_g5407 ( .A(I13937), .ZN(g5407) );
INV_X32 U_I13940 ( .A(g1739), .ZN(I13940) );
INV_X32 U_g5408 ( .A(I13940), .ZN(g5408) );
INV_X32 U_I13943 ( .A(g2418), .ZN(I13943) );
INV_X32 U_g5409 ( .A(I13943), .ZN(g5409) );
INV_X32 U_g5410 ( .A(g3079), .ZN(g5410) );
INV_X32 U_I13947 ( .A(g391), .ZN(I13947) );
INV_X32 U_g5411 ( .A(I13947), .ZN(g5411) );
INV_X32 U_I13950 ( .A(g1063), .ZN(I13950) );
INV_X32 U_g5412 ( .A(I13950), .ZN(g5412) );
INV_X32 U_I13953 ( .A(g1075), .ZN(I13953) );
INV_X32 U_g5413 ( .A(I13953), .ZN(g5413) );
INV_X32 U_I13956 ( .A(g1742), .ZN(I13956) );
INV_X32 U_g5414 ( .A(I13956), .ZN(g5414) );
INV_X32 U_I13959 ( .A(g1754), .ZN(I13959) );
INV_X32 U_g5415 ( .A(I13959), .ZN(g5415) );
INV_X32 U_I13962 ( .A(g2421), .ZN(I13962) );
INV_X32 U_g5416 ( .A(I13962), .ZN(g5416) );
INV_X32 U_I13965 ( .A(g2433), .ZN(I13965) );
INV_X32 U_g5417 ( .A(I13965), .ZN(g5417) );
INV_X32 U_I13968 ( .A(g1078), .ZN(I13968) );
INV_X32 U_g5418 ( .A(I13968), .ZN(g5418) );
INV_X32 U_I13971 ( .A(g1757), .ZN(I13971) );
INV_X32 U_g5419 ( .A(I13971), .ZN(g5419) );
INV_X32 U_I13974 ( .A(g1769), .ZN(I13974) );
INV_X32 U_g5420 ( .A(I13974), .ZN(g5420) );
INV_X32 U_I13977 ( .A(g2436), .ZN(I13977) );
INV_X32 U_g5421 ( .A(I13977), .ZN(g5421) );
INV_X32 U_I13980 ( .A(g2448), .ZN(I13980) );
INV_X32 U_g5422 ( .A(I13980), .ZN(g5422) );
INV_X32 U_g5423 ( .A(g2879), .ZN(g5423) );
INV_X32 U_I13984 ( .A(g1772), .ZN(I13984) );
INV_X32 U_g5424 ( .A(I13984), .ZN(g5424) );
INV_X32 U_I13987 ( .A(g2451), .ZN(I13987) );
INV_X32 U_g5425 ( .A(I13987), .ZN(g5425) );
INV_X32 U_I13990 ( .A(g2463), .ZN(I13990) );
INV_X32 U_g5426 ( .A(I13990), .ZN(g5426) );
INV_X32 U_I13993 ( .A(g2466), .ZN(I13993) );
INV_X32 U_g5427 ( .A(I13993), .ZN(g5427) );
INV_X32 U_g5428 ( .A(g3210), .ZN(g5428) );
INV_X32 U_g5431 ( .A(g3211), .ZN(g5431) );
INV_X32 U_g5434 ( .A(g3084), .ZN(g5434) );
INV_X32 U_I13999 ( .A(g276), .ZN(I13999) );
INV_X32 U_g5437 ( .A(I13999), .ZN(g5437) );
INV_X32 U_I14002 ( .A(g276), .ZN(I14002) );
INV_X32 U_g5438 ( .A(I14002), .ZN(g5438) );
INV_X32 U_g5469 ( .A(g3085), .ZN(g5469) );
INV_X32 U_I14006 ( .A(g963), .ZN(I14006) );
INV_X32 U_g5472 ( .A(I14006), .ZN(g5472) );
INV_X32 U_I14009 ( .A(g963), .ZN(I14009) );
INV_X32 U_g5473 ( .A(I14009), .ZN(g5473) );
INV_X32 U_g5504 ( .A(g3086), .ZN(g5504) );
INV_X32 U_g5507 ( .A(g3155), .ZN(g5507) );
INV_X32 U_I14014 ( .A(g499), .ZN(I14014) );
INV_X32 U_g5508 ( .A(I14014), .ZN(g5508) );
INV_X32 U_I14017 ( .A(g1657), .ZN(I14017) );
INV_X32 U_g5511 ( .A(I14017), .ZN(g5511) );
INV_X32 U_I14020 ( .A(g1657), .ZN(I14020) );
INV_X32 U_g5512 ( .A(I14020), .ZN(g5512) );
INV_X32 U_g5543 ( .A(g3087), .ZN(g5543) );
INV_X32 U_g5546 ( .A(g3164), .ZN(g5546) );
INV_X32 U_g5547 ( .A(g101), .ZN(g5547) );
INV_X32 U_g5548 ( .A(g105), .ZN(g5548) );
INV_X32 U_I14027 ( .A(g182), .ZN(I14027) );
INV_X32 U_g5549 ( .A(I14027), .ZN(g5549) );
INV_X32 U_I14030 ( .A(g182), .ZN(I14030) );
INV_X32 U_g5550 ( .A(I14030), .ZN(g5550) );
INV_X32 U_g5551 ( .A(g514), .ZN(g5551) );
INV_X32 U_I14034 ( .A(g1186), .ZN(I14034) );
INV_X32 U_g5552 ( .A(I14034), .ZN(g5552) );
INV_X32 U_I14037 ( .A(g2351), .ZN(I14037) );
INV_X32 U_g5555 ( .A(I14037), .ZN(g5555) );
INV_X32 U_I14040 ( .A(g2351), .ZN(I14040) );
INV_X32 U_g5556 ( .A(I14040), .ZN(g5556) );
INV_X32 U_g5587 ( .A(g3091), .ZN(g5587) );
INV_X32 U_g5590 ( .A(g3158), .ZN(g5590) );
INV_X32 U_g5591 ( .A(g3173), .ZN(g5591) );
INV_X32 U_g5592 ( .A(g515), .ZN(g5592) );
INV_X32 U_g5593 ( .A(g789), .ZN(g5593) );
INV_X32 U_g5594 ( .A(g793), .ZN(g5594) );
INV_X32 U_I14049 ( .A(g870), .ZN(I14049) );
INV_X32 U_g5595 ( .A(I14049), .ZN(g5595) );
INV_X32 U_I14052 ( .A(g870), .ZN(I14052) );
INV_X32 U_g5596 ( .A(I14052), .ZN(g5596) );
INV_X32 U_g5597 ( .A(g1200), .ZN(g5597) );
INV_X32 U_I14056 ( .A(g1880), .ZN(I14056) );
INV_X32 U_g5598 ( .A(I14056), .ZN(g5598) );
INV_X32 U_g5601 ( .A(g3092), .ZN(g5601) );
INV_X32 U_g5604 ( .A(g3167), .ZN(g5604) );
INV_X32 U_g5605 ( .A(g3182), .ZN(g5605) );
INV_X32 U_g5606 ( .A(g79), .ZN(g5606) );
INV_X32 U_g5609 ( .A(g1201), .ZN(g5609) );
INV_X32 U_g5610 ( .A(g1476), .ZN(g5610) );
INV_X32 U_g5611 ( .A(g1481), .ZN(g5611) );
INV_X32 U_I14066 ( .A(g1564), .ZN(I14066) );
INV_X32 U_g5612 ( .A(I14066), .ZN(g5612) );
INV_X32 U_I14069 ( .A(g1564), .ZN(I14069) );
INV_X32 U_g5613 ( .A(I14069), .ZN(g5613) );
INV_X32 U_g5614 ( .A(g1894), .ZN(g5614) );
INV_X32 U_I14073 ( .A(g2574), .ZN(I14073) );
INV_X32 U_g5615 ( .A(I14073), .ZN(g5615) );
INV_X32 U_g5618 ( .A(g3093), .ZN(g5618) );
INV_X32 U_g5621 ( .A(g3161), .ZN(g5621) );
INV_X32 U_g5622 ( .A(g3176), .ZN(g5622) );
INV_X32 U_g5623 ( .A(g70), .ZN(g5623) );
INV_X32 U_g5626 ( .A(g121), .ZN(g5626) );
INV_X32 U_g5627 ( .A(g125), .ZN(g5627) );
INV_X32 U_g5628 ( .A(g300), .ZN(g5628) );
INV_X32 U_I14083 ( .A(g325), .ZN(I14083) );
INV_X32 U_g5629 ( .A(I14083), .ZN(g5629) );
INV_X32 U_g5631 ( .A(g767), .ZN(g5631) );
INV_X32 U_g5634 ( .A(g1895), .ZN(g5634) );
INV_X32 U_g5635 ( .A(g2170), .ZN(g5635) );
INV_X32 U_g5636 ( .A(g2175), .ZN(g5636) );
INV_X32 U_I14091 ( .A(g2258), .ZN(I14091) );
INV_X32 U_g5637 ( .A(I14091), .ZN(g5637) );
INV_X32 U_I14094 ( .A(g2258), .ZN(I14094) );
INV_X32 U_g5638 ( .A(I14094), .ZN(g5638) );
INV_X32 U_g5639 ( .A(g2588), .ZN(g5639) );
INV_X32 U_g5640 ( .A(g3170), .ZN(g5640) );
INV_X32 U_g5641 ( .A(g3185), .ZN(g5641) );
INV_X32 U_g5642 ( .A(g61), .ZN(g5642) );
INV_X32 U_g5645 ( .A(g101), .ZN(g5645) );
INV_X32 U_g5646 ( .A(g213), .ZN(g5646) );
INV_X32 U_g5647 ( .A(g301), .ZN(g5647) );
INV_X32 U_I14104 ( .A(g331), .ZN(I14104) );
INV_X32 U_g5648 ( .A(I14104), .ZN(g5648) );
INV_X32 U_g5651 ( .A(g758), .ZN(g5651) );
INV_X32 U_g5654 ( .A(g809), .ZN(g5654) );
INV_X32 U_g5655 ( .A(g813), .ZN(g5655) );
INV_X32 U_g5656 ( .A(g987), .ZN(g5656) );
INV_X32 U_I14113 ( .A(g1012), .ZN(I14113) );
INV_X32 U_g5657 ( .A(I14113), .ZN(g5657) );
INV_X32 U_g5659 ( .A(g1453), .ZN(g5659) );
INV_X32 U_g5662 ( .A(g2589), .ZN(g5662) );
INV_X32 U_g5663 ( .A(g3179), .ZN(g5663) );
INV_X32 U_g5664 ( .A(g65), .ZN(g5664) );
INV_X32 U_g5665 ( .A(g105), .ZN(g5665) );
INV_X32 U_g5666 ( .A(g216), .ZN(g5666) );
INV_X32 U_g5667 ( .A(g222), .ZN(g5667) );
INV_X32 U_g5668 ( .A(g299), .ZN(g5668) );
INV_X32 U_g5675 ( .A(g302), .ZN(g5675) );
INV_X32 U_g5679 ( .A(g506), .ZN(g5679) );
INV_X32 U_g5680 ( .A(g749), .ZN(g5680) );
INV_X32 U_g5683 ( .A(g789), .ZN(g5683) );
INV_X32 U_g5684 ( .A(g900), .ZN(g5684) );
INV_X32 U_g5685 ( .A(g988), .ZN(g5685) );
INV_X32 U_I14134 ( .A(g1018), .ZN(I14134) );
INV_X32 U_g5686 ( .A(I14134), .ZN(g5686) );
INV_X32 U_g5689 ( .A(g1444), .ZN(g5689) );
INV_X32 U_g5692 ( .A(g1501), .ZN(g5692) );
INV_X32 U_g5693 ( .A(g1506), .ZN(g5693) );
INV_X32 U_g5694 ( .A(g1681), .ZN(g5694) );
INV_X32 U_I14143 ( .A(g1706), .ZN(I14143) );
INV_X32 U_g5695 ( .A(I14143), .ZN(g5695) );
INV_X32 U_g5697 ( .A(g2147), .ZN(g5697) );
INV_X32 U_g5700 ( .A(g3088), .ZN(g5700) );
INV_X32 U_I14149 ( .A(g3231), .ZN(I14149) );
INV_X32 U_g5701 ( .A(I14149), .ZN(g5701) );
INV_X32 U_g5702 ( .A(g56), .ZN(g5702) );
INV_X32 U_g5703 ( .A(g109), .ZN(g5703) );
INV_X32 U_g5704 ( .A(g219), .ZN(g5704) );
INV_X32 U_g5705 ( .A(g225), .ZN(g5705) );
INV_X32 U_g5706 ( .A(g231), .ZN(g5706) );
INV_X32 U_g5707 ( .A(g109), .ZN(g5707) );
INV_X32 U_g5708 ( .A(g303), .ZN(g5708) );
INV_X32 U_g5712 ( .A(g305), .ZN(g5712) );
INV_X32 U_I14163 ( .A(g113), .ZN(I14163) );
INV_X32 U_g5713 ( .A(I14163), .ZN(g5713) );
INV_X32 U_g5714 ( .A(g507), .ZN(g5714) );
INV_X32 U_g5715 ( .A(g541), .ZN(g5715) );
INV_X32 U_g5716 ( .A(g753), .ZN(g5716) );
INV_X32 U_g5717 ( .A(g793), .ZN(g5717) );
INV_X32 U_g5718 ( .A(g903), .ZN(g5718) );
INV_X32 U_g5719 ( .A(g909), .ZN(g5719) );
INV_X32 U_g5720 ( .A(g986), .ZN(g5720) );
INV_X32 U_g5727 ( .A(g989), .ZN(g5727) );
INV_X32 U_g5731 ( .A(g1192), .ZN(g5731) );
INV_X32 U_g5732 ( .A(g1435), .ZN(g5732) );
INV_X32 U_g5735 ( .A(g1476), .ZN(g5735) );
INV_X32 U_g5736 ( .A(g1594), .ZN(g5736) );
INV_X32 U_g5737 ( .A(g1682), .ZN(g5737) );
INV_X32 U_I14182 ( .A(g1712), .ZN(I14182) );
INV_X32 U_g5738 ( .A(I14182), .ZN(g5738) );
INV_X32 U_g5741 ( .A(g2138), .ZN(g5741) );
INV_X32 U_g5744 ( .A(g2195), .ZN(g5744) );
INV_X32 U_g5745 ( .A(g2200), .ZN(g5745) );
INV_X32 U_g5746 ( .A(g2375), .ZN(g5746) );
INV_X32 U_I14191 ( .A(g2400), .ZN(I14191) );
INV_X32 U_g5747 ( .A(I14191), .ZN(g5747) );
INV_X32 U_I14195 ( .A(g3212), .ZN(I14195) );
INV_X32 U_g5749 ( .A(I14195), .ZN(g5749) );
INV_X32 U_g5750 ( .A(g92), .ZN(g5750) );
INV_X32 U_g5751 ( .A(g52), .ZN(g5751) );
INV_X32 U_g5752 ( .A(g113), .ZN(g5752) );
INV_X32 U_g5753 ( .A(g228), .ZN(g5753) );
INV_X32 U_g5754 ( .A(g234), .ZN(g5754) );
INV_X32 U_g5755 ( .A(g240), .ZN(g5755) );
INV_X32 U_g5756 ( .A(g304), .ZN(g5756) );
INV_X32 U_g5759 ( .A(g508), .ZN(g5759) );
INV_X32 U_g5760 ( .A(g744), .ZN(g5760) );
INV_X32 U_g5761 ( .A(g797), .ZN(g5761) );
INV_X32 U_g5762 ( .A(g906), .ZN(g5762) );
INV_X32 U_g5763 ( .A(g912), .ZN(g5763) );
INV_X32 U_g5764 ( .A(g918), .ZN(g5764) );
INV_X32 U_g5765 ( .A(g797), .ZN(g5765) );
INV_X32 U_g5766 ( .A(g990), .ZN(g5766) );
INV_X32 U_g5770 ( .A(g992), .ZN(g5770) );
INV_X32 U_I14219 ( .A(g801), .ZN(I14219) );
INV_X32 U_g5771 ( .A(I14219), .ZN(g5771) );
INV_X32 U_g5772 ( .A(g1193), .ZN(g5772) );
INV_X32 U_g5773 ( .A(g1227), .ZN(g5773) );
INV_X32 U_g5774 ( .A(g1439), .ZN(g5774) );
INV_X32 U_g5775 ( .A(g1481), .ZN(g5775) );
INV_X32 U_g5776 ( .A(g1597), .ZN(g5776) );
INV_X32 U_g5777 ( .A(g1603), .ZN(g5777) );
INV_X32 U_g5778 ( .A(g1680), .ZN(g5778) );
INV_X32 U_g5785 ( .A(g1683), .ZN(g5785) );
INV_X32 U_g5789 ( .A(g1886), .ZN(g5789) );
INV_X32 U_g5790 ( .A(g2129), .ZN(g5790) );
INV_X32 U_g5793 ( .A(g2170), .ZN(g5793) );
INV_X32 U_g5794 ( .A(g2288), .ZN(g5794) );
INV_X32 U_g5795 ( .A(g2376), .ZN(g5795) );
INV_X32 U_I14238 ( .A(g2406), .ZN(I14238) );
INV_X32 U_g5796 ( .A(I14238), .ZN(g5796) );
INV_X32 U_I14243 ( .A(g3221), .ZN(I14243) );
INV_X32 U_g5799 ( .A(I14243), .ZN(g5799) );
INV_X32 U_I14246 ( .A(g3227), .ZN(I14246) );
INV_X32 U_g5800 ( .A(I14246), .ZN(g5800) );
INV_X32 U_I14249 ( .A(g3216), .ZN(I14249) );
INV_X32 U_g5801 ( .A(I14249), .ZN(g5801) );
INV_X32 U_g5802 ( .A(g83), .ZN(g5802) );
INV_X32 U_g5803 ( .A(g117), .ZN(g5803) );
INV_X32 U_g5804 ( .A(g237), .ZN(g5804) );
INV_X32 U_g5805 ( .A(g243), .ZN(g5805) );
INV_X32 U_g5806 ( .A(g249), .ZN(g5806) );
INV_X32 U_g5808 ( .A(g509), .ZN(g5808) );
INV_X32 U_g5809 ( .A(g780), .ZN(g5809) );
INV_X32 U_g5810 ( .A(g740), .ZN(g5810) );
INV_X32 U_g5811 ( .A(g801), .ZN(g5811) );
INV_X32 U_g5812 ( .A(g915), .ZN(g5812) );
INV_X32 U_g5813 ( .A(g921), .ZN(g5813) );
INV_X32 U_g5814 ( .A(g927), .ZN(g5814) );
INV_X32 U_g5815 ( .A(g991), .ZN(g5815) );
INV_X32 U_g5818 ( .A(g1194), .ZN(g5818) );
INV_X32 U_g5819 ( .A(g1430), .ZN(g5819) );
INV_X32 U_g5820 ( .A(g1486), .ZN(g5820) );
INV_X32 U_g5821 ( .A(g1600), .ZN(g5821) );
INV_X32 U_g5822 ( .A(g1606), .ZN(g5822) );
INV_X32 U_g5823 ( .A(g1612), .ZN(g5823) );
INV_X32 U_g5824 ( .A(g1486), .ZN(g5824) );
INV_X32 U_g5825 ( .A(g1684), .ZN(g5825) );
INV_X32 U_g5829 ( .A(g1686), .ZN(g5829) );
INV_X32 U_I14280 ( .A(g1491), .ZN(I14280) );
INV_X32 U_g5830 ( .A(I14280), .ZN(g5830) );
INV_X32 U_g5831 ( .A(g1887), .ZN(g5831) );
INV_X32 U_g5832 ( .A(g1921), .ZN(g5832) );
INV_X32 U_g5833 ( .A(g2133), .ZN(g5833) );
INV_X32 U_g5834 ( .A(g2175), .ZN(g5834) );
INV_X32 U_g5835 ( .A(g2291), .ZN(g5835) );
INV_X32 U_g5836 ( .A(g2297), .ZN(g5836) );
INV_X32 U_g5837 ( .A(g2374), .ZN(g5837) );
INV_X32 U_g5844 ( .A(g2377), .ZN(g5844) );
INV_X32 U_g5848 ( .A(g2580), .ZN(g5848) );
INV_X32 U_I14295 ( .A(g3228), .ZN(I14295) );
INV_X32 U_g5849 ( .A(I14295), .ZN(g5849) );
INV_X32 U_I14298 ( .A(g3217), .ZN(I14298) );
INV_X32 U_g5850 ( .A(I14298), .ZN(g5850) );
INV_X32 U_g5851 ( .A(g74), .ZN(g5851) );
INV_X32 U_g5852 ( .A(g121), .ZN(g5852) );
INV_X32 U_g5853 ( .A(g246), .ZN(g5853) );
INV_X32 U_g5854 ( .A(g252), .ZN(g5854) );
INV_X32 U_g5855 ( .A(g258), .ZN(g5855) );
INV_X32 U_I14306 ( .A(g97), .ZN(I14306) );
INV_X32 U_g5856 ( .A(I14306), .ZN(g5856) );
INV_X32 U_g5857 ( .A(g538), .ZN(g5857) );
INV_X32 U_g5858 ( .A(g771), .ZN(g5858) );
INV_X32 U_g5859 ( .A(g805), .ZN(g5859) );
INV_X32 U_g5860 ( .A(g924), .ZN(g5860) );
INV_X32 U_g5861 ( .A(g930), .ZN(g5861) );
INV_X32 U_g5862 ( .A(g936), .ZN(g5862) );
INV_X32 U_g5864 ( .A(g1195), .ZN(g5864) );
INV_X32 U_g5865 ( .A(g1466), .ZN(g5865) );
INV_X32 U_g5866 ( .A(g1426), .ZN(g5866) );
INV_X32 U_g5867 ( .A(g1491), .ZN(g5867) );
INV_X32 U_g5868 ( .A(g1609), .ZN(g5868) );
INV_X32 U_g5869 ( .A(g1615), .ZN(g5869) );
INV_X32 U_g5870 ( .A(g1621), .ZN(g5870) );
INV_X32 U_g5871 ( .A(g1685), .ZN(g5871) );
INV_X32 U_g5874 ( .A(g1888), .ZN(g5874) );
INV_X32 U_g5875 ( .A(g2124), .ZN(g5875) );
INV_X32 U_g5876 ( .A(g2180), .ZN(g5876) );
INV_X32 U_g5877 ( .A(g2294), .ZN(g5877) );
INV_X32 U_g5878 ( .A(g2300), .ZN(g5878) );
INV_X32 U_g5879 ( .A(g2306), .ZN(g5879) );
INV_X32 U_g5880 ( .A(g2180), .ZN(g5880) );
INV_X32 U_g5881 ( .A(g2378), .ZN(g5881) );
INV_X32 U_g5885 ( .A(g2380), .ZN(g5885) );
INV_X32 U_I14338 ( .A(g2185), .ZN(I14338) );
INV_X32 U_g5886 ( .A(I14338), .ZN(g5886) );
INV_X32 U_g5887 ( .A(g2581), .ZN(g5887) );
INV_X32 U_g5888 ( .A(g2615), .ZN(g5888) );
INV_X32 U_I14343 ( .A(g3219), .ZN(I14343) );
INV_X32 U_g5889 ( .A(I14343), .ZN(g5889) );
INV_X32 U_g5890 ( .A(g88), .ZN(g5890) );
INV_X32 U_g5893 ( .A(g125), .ZN(g5893) );
INV_X32 U_g5894 ( .A(g186), .ZN(g5894) );
INV_X32 U_g5895 ( .A(g255), .ZN(g5895) );
INV_X32 U_g5896 ( .A(g261), .ZN(g5896) );
INV_X32 U_g5897 ( .A(g267), .ZN(g5897) );
INV_X32 U_g5898 ( .A(g762), .ZN(g5898) );
INV_X32 U_g5899 ( .A(g809), .ZN(g5899) );
INV_X32 U_g5900 ( .A(g933), .ZN(g5900) );
INV_X32 U_g5901 ( .A(g939), .ZN(g5901) );
INV_X32 U_g5902 ( .A(g945), .ZN(g5902) );
INV_X32 U_I14357 ( .A(g785), .ZN(I14357) );
INV_X32 U_g5903 ( .A(I14357), .ZN(g5903) );
INV_X32 U_g5904 ( .A(g1224), .ZN(g5904) );
INV_X32 U_g5905 ( .A(g1457), .ZN(g5905) );
INV_X32 U_g5906 ( .A(g1496), .ZN(g5906) );
INV_X32 U_g5907 ( .A(g1618), .ZN(g5907) );
INV_X32 U_g5908 ( .A(g1624), .ZN(g5908) );
INV_X32 U_g5909 ( .A(g1630), .ZN(g5909) );
INV_X32 U_g5911 ( .A(g1889), .ZN(g5911) );
INV_X32 U_g5912 ( .A(g2160), .ZN(g5912) );
INV_X32 U_g5913 ( .A(g2120), .ZN(g5913) );
INV_X32 U_g5914 ( .A(g2185), .ZN(g5914) );
INV_X32 U_g5915 ( .A(g2303), .ZN(g5915) );
INV_X32 U_g5916 ( .A(g2309), .ZN(g5916) );
INV_X32 U_g5917 ( .A(g2315), .ZN(g5917) );
INV_X32 U_g5918 ( .A(g2379), .ZN(g5918) );
INV_X32 U_g5921 ( .A(g2582), .ZN(g5921) );
INV_X32 U_I14378 ( .A(g3234), .ZN(I14378) );
INV_X32 U_g5922 ( .A(I14378), .ZN(g5922) );
INV_X32 U_I14381 ( .A(g3223), .ZN(I14381) );
INV_X32 U_g5923 ( .A(I14381), .ZN(g5923) );
INV_X32 U_I14384 ( .A(g3218), .ZN(I14384) );
INV_X32 U_g5924 ( .A(I14384), .ZN(g5924) );
INV_X32 U_g5925 ( .A(g189), .ZN(g5925) );
INV_X32 U_g5926 ( .A(g195), .ZN(g5926) );
INV_X32 U_g5927 ( .A(g264), .ZN(g5927) );
INV_X32 U_g5928 ( .A(g270), .ZN(g5928) );
INV_X32 U_g5929 ( .A(g776), .ZN(g5929) );
INV_X32 U_g5932 ( .A(g813), .ZN(g5932) );
INV_X32 U_g5933 ( .A(g873), .ZN(g5933) );
INV_X32 U_g5934 ( .A(g942), .ZN(g5934) );
INV_X32 U_g5935 ( .A(g948), .ZN(g5935) );
INV_X32 U_g5936 ( .A(g954), .ZN(g5936) );
INV_X32 U_g5937 ( .A(g1448), .ZN(g5937) );
INV_X32 U_g5938 ( .A(g1501), .ZN(g5938) );
INV_X32 U_g5939 ( .A(g1627), .ZN(g5939) );
INV_X32 U_g5940 ( .A(g1633), .ZN(g5940) );
INV_X32 U_g5941 ( .A(g1639), .ZN(g5941) );
INV_X32 U_I14402 ( .A(g1471), .ZN(I14402) );
INV_X32 U_g5942 ( .A(I14402), .ZN(g5942) );
INV_X32 U_g5943 ( .A(g1918), .ZN(g5943) );
INV_X32 U_g5944 ( .A(g2151), .ZN(g5944) );
INV_X32 U_g5945 ( .A(g2190), .ZN(g5945) );
INV_X32 U_g5946 ( .A(g2312), .ZN(g5946) );
INV_X32 U_g5947 ( .A(g2318), .ZN(g5947) );
INV_X32 U_g5948 ( .A(g2324), .ZN(g5948) );
INV_X32 U_g5950 ( .A(g2583), .ZN(g5950) );
INV_X32 U_I14413 ( .A(g3233), .ZN(I14413) );
INV_X32 U_g5951 ( .A(I14413), .ZN(g5951) );
INV_X32 U_I14416 ( .A(g3222), .ZN(I14416) );
INV_X32 U_g5952 ( .A(I14416), .ZN(g5952) );
INV_X32 U_g5953 ( .A(g97), .ZN(g5953) );
INV_X32 U_g5954 ( .A(g192), .ZN(g5954) );
INV_X32 U_g5955 ( .A(g198), .ZN(g5955) );
INV_X32 U_g5956 ( .A(g204), .ZN(g5956) );
INV_X32 U_g5957 ( .A(g273), .ZN(g5957) );
INV_X32 U_I14424 ( .A(g117), .ZN(I14424) );
INV_X32 U_g5958 ( .A(I14424), .ZN(g5958) );
INV_X32 U_g5959 ( .A(g876), .ZN(g5959) );
INV_X32 U_g5960 ( .A(g882), .ZN(g5960) );
INV_X32 U_g5961 ( .A(g951), .ZN(g5961) );
INV_X32 U_g5962 ( .A(g957), .ZN(g5962) );
INV_X32 U_g5963 ( .A(g1462), .ZN(g5963) );
INV_X32 U_g5966 ( .A(g1506), .ZN(g5966) );
INV_X32 U_g5967 ( .A(g1567), .ZN(g5967) );
INV_X32 U_g5968 ( .A(g1636), .ZN(g5968) );
INV_X32 U_g5969 ( .A(g1642), .ZN(g5969) );
INV_X32 U_g5970 ( .A(g1648), .ZN(g5970) );
INV_X32 U_g5971 ( .A(g2142), .ZN(g5971) );
INV_X32 U_g5972 ( .A(g2195), .ZN(g5972) );
INV_X32 U_g5973 ( .A(g2321), .ZN(g5973) );
INV_X32 U_g5974 ( .A(g2327), .ZN(g5974) );
INV_X32 U_g5975 ( .A(g2333), .ZN(g5975) );
INV_X32 U_I14442 ( .A(g2165), .ZN(I14442) );
INV_X32 U_g5976 ( .A(I14442), .ZN(g5976) );
INV_X32 U_g5977 ( .A(g2612), .ZN(g5977) );
INV_X32 U_I14446 ( .A(g3230), .ZN(I14446) );
INV_X32 U_g5978 ( .A(I14446), .ZN(g5978) );
INV_X32 U_I14449 ( .A(g3224), .ZN(I14449) );
INV_X32 U_g5979 ( .A(I14449), .ZN(g5979) );
INV_X32 U_g5980 ( .A(g201), .ZN(g5980) );
INV_X32 U_g5981 ( .A(g207), .ZN(g5981) );
INV_X32 U_g5982 ( .A(g785), .ZN(g5982) );
INV_X32 U_g5983 ( .A(g879), .ZN(g5983) );
INV_X32 U_g5984 ( .A(g885), .ZN(g5984) );
INV_X32 U_g5985 ( .A(g891), .ZN(g5985) );
INV_X32 U_g5986 ( .A(g960), .ZN(g5986) );
INV_X32 U_I14459 ( .A(g805), .ZN(I14459) );
INV_X32 U_g5987 ( .A(I14459), .ZN(g5987) );
INV_X32 U_g5988 ( .A(g1570), .ZN(g5988) );
INV_X32 U_g5989 ( .A(g1576), .ZN(g5989) );
INV_X32 U_g5990 ( .A(g1645), .ZN(g5990) );
INV_X32 U_g5991 ( .A(g1651), .ZN(g5991) );
INV_X32 U_g5992 ( .A(g2156), .ZN(g5992) );
INV_X32 U_g5995 ( .A(g2200), .ZN(g5995) );
INV_X32 U_g5996 ( .A(g2261), .ZN(g5996) );
INV_X32 U_g5997 ( .A(g2330), .ZN(g5997) );
INV_X32 U_g5998 ( .A(g2336), .ZN(g5998) );
INV_X32 U_g5999 ( .A(g2342), .ZN(g5999) );
INV_X32 U_I14472 ( .A(g3080), .ZN(I14472) );
INV_X32 U_g6000 ( .A(I14472), .ZN(g6000) );
INV_X32 U_I14475 ( .A(g3225), .ZN(I14475) );
INV_X32 U_g6014 ( .A(I14475), .ZN(g6014) );
INV_X32 U_I14478 ( .A(g3213), .ZN(I14478) );
INV_X32 U_g6015 ( .A(I14478), .ZN(g6015) );
INV_X32 U_g6016 ( .A(g210), .ZN(g6016) );
INV_X32 U_g6017 ( .A(g888), .ZN(g6017) );
INV_X32 U_g6018 ( .A(g894), .ZN(g6018) );
INV_X32 U_g6019 ( .A(g1471), .ZN(g6019) );
INV_X32 U_g6020 ( .A(g1573), .ZN(g6020) );
INV_X32 U_g6021 ( .A(g1579), .ZN(g6021) );
INV_X32 U_g6022 ( .A(g1585), .ZN(g6022) );
INV_X32 U_g6023 ( .A(g1654), .ZN(g6023) );
INV_X32 U_I14489 ( .A(g1496), .ZN(I14489) );
INV_X32 U_g6024 ( .A(I14489), .ZN(g6024) );
INV_X32 U_g6025 ( .A(g2264), .ZN(g6025) );
INV_X32 U_g6026 ( .A(g2270), .ZN(g6026) );
INV_X32 U_g6027 ( .A(g2339), .ZN(g6027) );
INV_X32 U_g6028 ( .A(g2345), .ZN(g6028) );
INV_X32 U_I14496 ( .A(g3226), .ZN(I14496) );
INV_X32 U_g6029 ( .A(I14496), .ZN(g6029) );
INV_X32 U_I14499 ( .A(g3214), .ZN(I14499) );
INV_X32 U_g6030 ( .A(I14499), .ZN(g6030) );
INV_X32 U_I14502 ( .A(g471), .ZN(I14502) );
INV_X32 U_g6031 ( .A(I14502), .ZN(g6031) );
INV_X32 U_g6032 ( .A(g897), .ZN(g6032) );
INV_X32 U_g6033 ( .A(g1582), .ZN(g6033) );
INV_X32 U_g6034 ( .A(g1588), .ZN(g6034) );
INV_X32 U_g6035 ( .A(g2165), .ZN(g6035) );
INV_X32 U_g6036 ( .A(g2267), .ZN(g6036) );
INV_X32 U_g6037 ( .A(g2273), .ZN(g6037) );
INV_X32 U_g6038 ( .A(g2279), .ZN(g6038) );
INV_X32 U_g6039 ( .A(g2348), .ZN(g6039) );
INV_X32 U_I14513 ( .A(g2190), .ZN(I14513) );
INV_X32 U_g6040 ( .A(I14513), .ZN(g6040) );
INV_X32 U_I14516 ( .A(g3215), .ZN(I14516) );
INV_X32 U_g6041 ( .A(I14516), .ZN(g6041) );
INV_X32 U_I14519 ( .A(g1158), .ZN(I14519) );
INV_X32 U_g6042 ( .A(I14519), .ZN(g6042) );
INV_X32 U_g6043 ( .A(g1591), .ZN(g6043) );
INV_X32 U_g6044 ( .A(g2276), .ZN(g6044) );
INV_X32 U_g6045 ( .A(g2282), .ZN(g6045) );
INV_X32 U_I14525 ( .A(g1852), .ZN(I14525) );
INV_X32 U_g6046 ( .A(I14525), .ZN(g6046) );
INV_X32 U_g6047 ( .A(g2285), .ZN(g6047) );
INV_X32 U_I14529 ( .A(g3142), .ZN(I14529) );
INV_X32 U_g6048 ( .A(I14529), .ZN(g6048) );
INV_X32 U_I14532 ( .A(g354), .ZN(I14532) );
INV_X32 U_g6051 ( .A(I14532), .ZN(g6051) );
INV_X32 U_I14535 ( .A(g2546), .ZN(I14535) );
INV_X32 U_g6052 ( .A(I14535), .ZN(g6052) );
INV_X32 U_I14538 ( .A(g369), .ZN(I14538) );
INV_X32 U_g6053 ( .A(I14538), .ZN(g6053) );
INV_X32 U_I14541 ( .A(g455), .ZN(I14541) );
INV_X32 U_g6054 ( .A(I14541), .ZN(g6054) );
INV_X32 U_I14544 ( .A(g1041), .ZN(I14544) );
INV_X32 U_g6055 ( .A(I14544), .ZN(g6055) );
INV_X32 U_I14547 ( .A(g384), .ZN(I14547) );
INV_X32 U_g6056 ( .A(I14547), .ZN(g6056) );
INV_X32 U_I14550 ( .A(g458), .ZN(I14550) );
INV_X32 U_g6057 ( .A(I14550), .ZN(g6057) );
INV_X32 U_I14553 ( .A(g1056), .ZN(I14553) );
INV_X32 U_g6058 ( .A(I14553), .ZN(g6058) );
INV_X32 U_I14556 ( .A(g1142), .ZN(I14556) );
INV_X32 U_g6059 ( .A(I14556), .ZN(g6059) );
INV_X32 U_I14559 ( .A(g1735), .ZN(I14559) );
INV_X32 U_g6060 ( .A(I14559), .ZN(g6060) );
INV_X32 U_I14562 ( .A(g398), .ZN(I14562) );
INV_X32 U_g6061 ( .A(I14562), .ZN(g6061) );
INV_X32 U_I14565 ( .A(g461), .ZN(I14565) );
INV_X32 U_g6062 ( .A(I14565), .ZN(g6062) );
INV_X32 U_I14568 ( .A(g1071), .ZN(I14568) );
INV_X32 U_g6063 ( .A(I14568), .ZN(g6063) );
INV_X32 U_I14571 ( .A(g1145), .ZN(I14571) );
INV_X32 U_g6064 ( .A(I14571), .ZN(g6064) );
INV_X32 U_I14574 ( .A(g1750), .ZN(I14574) );
INV_X32 U_g6065 ( .A(I14574), .ZN(g6065) );
INV_X32 U_I14577 ( .A(g1836), .ZN(I14577) );
INV_X32 U_g6066 ( .A(I14577), .ZN(g6066) );
INV_X32 U_I14580 ( .A(g2429), .ZN(I14580) );
INV_X32 U_g6067 ( .A(I14580), .ZN(g6067) );
INV_X32 U_g6068 ( .A(g499), .ZN(g6068) );
INV_X32 U_I14584 ( .A(g465), .ZN(I14584) );
INV_X32 U_g6079 ( .A(I14584), .ZN(g6079) );
INV_X32 U_I14587 ( .A(g1085), .ZN(I14587) );
INV_X32 U_g6080 ( .A(I14587), .ZN(g6080) );
INV_X32 U_I14590 ( .A(g1148), .ZN(I14590) );
INV_X32 U_g6081 ( .A(I14590), .ZN(g6081) );
INV_X32 U_I14593 ( .A(g1765), .ZN(I14593) );
INV_X32 U_g6082 ( .A(I14593), .ZN(g6082) );
INV_X32 U_I14596 ( .A(g1839), .ZN(I14596) );
INV_X32 U_g6083 ( .A(I14596), .ZN(g6083) );
INV_X32 U_I14599 ( .A(g2444), .ZN(I14599) );
INV_X32 U_g6084 ( .A(I14599), .ZN(g6084) );
INV_X32 U_I14602 ( .A(g2530), .ZN(I14602) );
INV_X32 U_g6085 ( .A(I14602), .ZN(g6085) );
INV_X32 U_I14605 ( .A(g468), .ZN(I14605) );
INV_X32 U_g6086 ( .A(I14605), .ZN(g6086) );
INV_X32 U_g6087 ( .A(g1186), .ZN(g6087) );
INV_X32 U_I14609 ( .A(g1152), .ZN(I14609) );
INV_X32 U_g6098 ( .A(I14609), .ZN(g6098) );
INV_X32 U_I14612 ( .A(g1779), .ZN(I14612) );
INV_X32 U_g6099 ( .A(I14612), .ZN(g6099) );
INV_X32 U_I14615 ( .A(g1842), .ZN(I14615) );
INV_X32 U_g6100 ( .A(I14615), .ZN(g6100) );
INV_X32 U_I14618 ( .A(g2459), .ZN(I14618) );
INV_X32 U_g6101 ( .A(I14618), .ZN(g6101) );
INV_X32 U_I14621 ( .A(g2533), .ZN(I14621) );
INV_X32 U_g6102 ( .A(I14621), .ZN(g6102) );
INV_X32 U_I14624 ( .A(g1155), .ZN(I14624) );
INV_X32 U_g6103 ( .A(I14624), .ZN(g6103) );
INV_X32 U_g6104 ( .A(g1880), .ZN(g6104) );
INV_X32 U_I14628 ( .A(g1846), .ZN(I14628) );
INV_X32 U_g6115 ( .A(I14628), .ZN(g6115) );
INV_X32 U_I14631 ( .A(g2473), .ZN(I14631) );
INV_X32 U_g6116 ( .A(I14631), .ZN(g6116) );
INV_X32 U_I14634 ( .A(g2536), .ZN(I14634) );
INV_X32 U_g6117 ( .A(I14634), .ZN(g6117) );
INV_X32 U_I14637 ( .A(g1849), .ZN(I14637) );
INV_X32 U_g6118 ( .A(I14637), .ZN(g6118) );
INV_X32 U_g6119 ( .A(g2574), .ZN(g6119) );
INV_X32 U_I14641 ( .A(g2540), .ZN(I14641) );
INV_X32 U_g6130 ( .A(I14641), .ZN(g6130) );
INV_X32 U_I14644 ( .A(g3142), .ZN(I14644) );
INV_X32 U_g6131 ( .A(I14644), .ZN(g6131) );
INV_X32 U_I14647 ( .A(g2543), .ZN(I14647) );
INV_X32 U_g6134 ( .A(I14647), .ZN(g6134) );
INV_X32 U_I14650 ( .A(g525), .ZN(I14650) );
INV_X32 U_g6135 ( .A(I14650), .ZN(g6135) );
INV_X32 U_g6136 ( .A(g672), .ZN(g6136) );
INV_X32 U_I14654 ( .A(g3220), .ZN(I14654) );
INV_X32 U_g6139 ( .A(I14654), .ZN(g6139) );
INV_X32 U_g6140 ( .A(g524), .ZN(g6140) );
INV_X32 U_g6141 ( .A(g554), .ZN(g6141) );
INV_X32 U_g6142 ( .A(g679), .ZN(g6142) );
INV_X32 U_I14660 ( .A(g1211), .ZN(I14660) );
INV_X32 U_g6145 ( .A(I14660), .ZN(g6145) );
INV_X32 U_g6146 ( .A(g1358), .ZN(g6146) );
INV_X32 U_g6149 ( .A(g3097), .ZN(g6149) );
INV_X32 U_I14665 ( .A(g3147), .ZN(I14665) );
INV_X32 U_g6153 ( .A(I14665), .ZN(g6153) );
INV_X32 U_I14668 ( .A(g3232), .ZN(I14668) );
INV_X32 U_g6156 ( .A(I14668), .ZN(g6156) );
INV_X32 U_g6157 ( .A(g686), .ZN(g6157) );
INV_X32 U_g6161 ( .A(g1210), .ZN(g6161) );
INV_X32 U_g6162 ( .A(g1240), .ZN(g6162) );
INV_X32 U_g6163 ( .A(g1365), .ZN(g6163) );
INV_X32 U_I14675 ( .A(g1905), .ZN(I14675) );
INV_X32 U_g6166 ( .A(I14675), .ZN(g6166) );
INV_X32 U_g6167 ( .A(g2052), .ZN(g6167) );
INV_X32 U_g6170 ( .A(g3098), .ZN(g6170) );
INV_X32 U_g6173 ( .A(g557), .ZN(g6173) );
INV_X32 U_g6177 ( .A(g633), .ZN(g6177) );
INV_X32 U_g6180 ( .A(g692), .ZN(g6180) );
INV_X32 U_g6183 ( .A(g291), .ZN(g6183) );
INV_X32 U_g6184 ( .A(g1372), .ZN(g6184) );
INV_X32 U_g6188 ( .A(g1904), .ZN(g6188) );
INV_X32 U_g6189 ( .A(g1934), .ZN(g6189) );
INV_X32 U_g6190 ( .A(g2059), .ZN(g6190) );
INV_X32 U_I14688 ( .A(g2599), .ZN(I14688) );
INV_X32 U_g6193 ( .A(I14688), .ZN(g6193) );
INV_X32 U_g6194 ( .A(g2746), .ZN(g6194) );
INV_X32 U_g6197 ( .A(g3099), .ZN(g6197) );
INV_X32 U_g6200 ( .A(g542), .ZN(g6200) );
INV_X32 U_g6201 ( .A(g646), .ZN(g6201) );
INV_X32 U_g6204 ( .A(g289), .ZN(g6204) );
INV_X32 U_g6205 ( .A(g1243), .ZN(g6205) );
INV_X32 U_g6209 ( .A(g1319), .ZN(g6209) );
INV_X32 U_g6212 ( .A(g1378), .ZN(g6212) );
INV_X32 U_g6215 ( .A(g978), .ZN(g6215) );
INV_X32 U_g6216 ( .A(g2066), .ZN(g6216) );
INV_X32 U_g6220 ( .A(g2598), .ZN(g6220) );
INV_X32 U_g6221 ( .A(g2628), .ZN(g6221) );
INV_X32 U_g6222 ( .A(g2753), .ZN(g6222) );
INV_X32 U_I14704 ( .A(g2818), .ZN(I14704) );
INV_X32 U_g6225 ( .A(I14704), .ZN(g6225) );
INV_X32 U_g6226 ( .A(g2818), .ZN(g6226) );
INV_X32 U_g6227 ( .A(g3100), .ZN(g6227) );
INV_X32 U_I14709 ( .A(g3229), .ZN(I14709) );
INV_X32 U_g6230 ( .A(I14709), .ZN(g6230) );
INV_X32 U_I14712 ( .A(g138), .ZN(I14712) );
INV_X32 U_g6231 ( .A(I14712), .ZN(g6231) );
INV_X32 U_I14715 ( .A(g138), .ZN(I14715) );
INV_X32 U_g6232 ( .A(I14715), .ZN(g6232) );
INV_X32 U_g6281 ( .A(g510), .ZN(g6281) );
INV_X32 U_g6284 ( .A(g640), .ZN(g6284) );
INV_X32 U_g6288 ( .A(g287), .ZN(g6288) );
INV_X32 U_g6289 ( .A(g1228), .ZN(g6289) );
INV_X32 U_g6290 ( .A(g1332), .ZN(g6290) );
INV_X32 U_g6293 ( .A(g976), .ZN(g6293) );
INV_X32 U_g6294 ( .A(g1937), .ZN(g6294) );
INV_X32 U_g6298 ( .A(g2013), .ZN(g6298) );
INV_X32 U_g6301 ( .A(g2072), .ZN(g6301) );
INV_X32 U_g6304 ( .A(g1672), .ZN(g6304) );
INV_X32 U_g6305 ( .A(g2760), .ZN(g6305) );
INV_X32 U_g6309 ( .A(g14), .ZN(g6309) );
INV_X32 U_g6310 ( .A(g3101), .ZN(g6310) );
INV_X32 U_I14731 ( .A(g135), .ZN(I14731) );
INV_X32 U_g6313 ( .A(I14731), .ZN(g6313) );
INV_X32 U_I14734 ( .A(g135), .ZN(I14734) );
INV_X32 U_g6314 ( .A(I14734), .ZN(g6314) );
INV_X32 U_g6363 ( .A(g653), .ZN(g6363) );
INV_X32 U_g6367 ( .A(g285), .ZN(g6367) );
INV_X32 U_I14739 ( .A(g826), .ZN(I14739) );
INV_X32 U_g6368 ( .A(I14739), .ZN(g6368) );
INV_X32 U_I14742 ( .A(g826), .ZN(I14742) );
INV_X32 U_g6369 ( .A(I14742), .ZN(g6369) );
INV_X32 U_g6418 ( .A(g1196), .ZN(g6418) );
INV_X32 U_g6421 ( .A(g1326), .ZN(g6421) );
INV_X32 U_g6425 ( .A(g974), .ZN(g6425) );
INV_X32 U_g6426 ( .A(g1922), .ZN(g6426) );
INV_X32 U_g6427 ( .A(g2026), .ZN(g6427) );
INV_X32 U_g6430 ( .A(g1670), .ZN(g6430) );
INV_X32 U_g6431 ( .A(g2631), .ZN(g6431) );
INV_X32 U_g6435 ( .A(g2707), .ZN(g6435) );
INV_X32 U_g6438 ( .A(g2766), .ZN(g6438) );
INV_X32 U_g6441 ( .A(g2366), .ZN(g6441) );
INV_X32 U_I14755 ( .A(g2821), .ZN(I14755) );
INV_X32 U_g6442 ( .A(I14755), .ZN(g6442) );
INV_X32 U_g6443 ( .A(g2821), .ZN(g6443) );
INV_X32 U_g6444 ( .A(g3102), .ZN(g6444) );
INV_X32 U_I14760 ( .A(g405), .ZN(I14760) );
INV_X32 U_g6447 ( .A(I14760), .ZN(g6447) );
INV_X32 U_I14763 ( .A(g405), .ZN(I14763) );
INV_X32 U_g6448 ( .A(I14763), .ZN(g6448) );
INV_X32 U_I14766 ( .A(g545), .ZN(I14766) );
INV_X32 U_g6485 ( .A(I14766), .ZN(g6485) );
INV_X32 U_I14769 ( .A(g545), .ZN(I14769) );
INV_X32 U_g6486 ( .A(I14769), .ZN(g6486) );
INV_X32 U_g6512 ( .A(g544), .ZN(g6512) );
INV_X32 U_g6513 ( .A(g660), .ZN(g6513) );
INV_X32 U_g6517 ( .A(g283), .ZN(g6517) );
INV_X32 U_I14775 ( .A(g823), .ZN(I14775) );
INV_X32 U_g6518 ( .A(I14775), .ZN(g6518) );
INV_X32 U_I14778 ( .A(g823), .ZN(I14778) );
INV_X32 U_g6519 ( .A(I14778), .ZN(g6519) );
INV_X32 U_g6568 ( .A(g1339), .ZN(g6568) );
INV_X32 U_g6572 ( .A(g972), .ZN(g6572) );
INV_X32 U_I14783 ( .A(g1520), .ZN(I14783) );
INV_X32 U_g6573 ( .A(I14783), .ZN(g6573) );
INV_X32 U_I14786 ( .A(g1520), .ZN(I14786) );
INV_X32 U_g6574 ( .A(I14786), .ZN(g6574) );
INV_X32 U_g6623 ( .A(g1890), .ZN(g6623) );
INV_X32 U_g6626 ( .A(g2020), .ZN(g6626) );
INV_X32 U_g6630 ( .A(g1668), .ZN(g6630) );
INV_X32 U_g6631 ( .A(g2616), .ZN(g6631) );
INV_X32 U_g6632 ( .A(g2720), .ZN(g6632) );
INV_X32 U_g6635 ( .A(g2364), .ZN(g6635) );
INV_X32 U_g6636 ( .A(g1491), .ZN(g6636) );
INV_X32 U_g6637 ( .A(g5), .ZN(g6637) );
INV_X32 U_g6638 ( .A(g3103), .ZN(g6638) );
INV_X32 U_g6641 ( .A(g113), .ZN(g6641) );
INV_X32 U_I14799 ( .A(g551), .ZN(I14799) );
INV_X32 U_g6642 ( .A(I14799), .ZN(g6642) );
INV_X32 U_I14802 ( .A(g551), .ZN(I14802) );
INV_X32 U_g6643 ( .A(I14802), .ZN(g6643) );
INV_X32 U_g6672 ( .A(g464), .ZN(g6672) );
INV_X32 U_g6675 ( .A(g458), .ZN(g6675) );
INV_X32 U_g6676 ( .A(g559), .ZN(g6676) );
INV_X32 U_I14808 ( .A(g623), .ZN(I14808) );
INV_X32 U_g6677 ( .A(I14808), .ZN(g6677) );
INV_X32 U_I14811 ( .A(g623), .ZN(I14811) );
INV_X32 U_g6678 ( .A(I14811), .ZN(g6678) );
INV_X32 U_g6707 ( .A(g666), .ZN(g6707) );
INV_X32 U_g6711 ( .A(g281), .ZN(g6711) );
INV_X32 U_I14816 ( .A(g1092), .ZN(I14816) );
INV_X32 U_g6712 ( .A(I14816), .ZN(g6712) );
INV_X32 U_I14819 ( .A(g1092), .ZN(I14819) );
INV_X32 U_g6713 ( .A(I14819), .ZN(g6713) );
INV_X32 U_I14822 ( .A(g1231), .ZN(I14822) );
INV_X32 U_g6750 ( .A(I14822), .ZN(g6750) );
INV_X32 U_I14825 ( .A(g1231), .ZN(I14825) );
INV_X32 U_g6751 ( .A(I14825), .ZN(g6751) );
INV_X32 U_g6776 ( .A(g1230), .ZN(g6776) );
INV_X32 U_g6777 ( .A(g1346), .ZN(g6777) );
INV_X32 U_g6781 ( .A(g970), .ZN(g6781) );
INV_X32 U_I14831 ( .A(g1517), .ZN(I14831) );
INV_X32 U_g6782 ( .A(I14831), .ZN(g6782) );
INV_X32 U_I14834 ( .A(g1517), .ZN(I14834) );
INV_X32 U_g6783 ( .A(I14834), .ZN(g6783) );
INV_X32 U_g6832 ( .A(g2033), .ZN(g6832) );
INV_X32 U_g6836 ( .A(g1666), .ZN(g6836) );
INV_X32 U_I14839 ( .A(g2214), .ZN(I14839) );
INV_X32 U_g6837 ( .A(I14839), .ZN(g6837) );
INV_X32 U_I14842 ( .A(g2214), .ZN(I14842) );
INV_X32 U_g6838 ( .A(I14842), .ZN(g6838) );
INV_X32 U_g6887 ( .A(g2584), .ZN(g6887) );
INV_X32 U_g6890 ( .A(g2714), .ZN(g6890) );
INV_X32 U_g6894 ( .A(g2362), .ZN(g6894) );
INV_X32 U_I14848 ( .A(g2824), .ZN(I14848) );
INV_X32 U_g6895 ( .A(I14848), .ZN(g6895) );
INV_X32 U_g6896 ( .A(g2824), .ZN(g6896) );
INV_X32 U_g6897 ( .A(g1486), .ZN(g6897) );
INV_X32 U_g6898 ( .A(g2993), .ZN(g6898) );
INV_X32 U_g6901 ( .A(g3006), .ZN(g6901) );
INV_X32 U_g6905 ( .A(g3104), .ZN(g6905) );
INV_X32 U_g6908 ( .A(g484), .ZN(g6908) );
INV_X32 U_I14857 ( .A(g626), .ZN(I14857) );
INV_X32 U_g6911 ( .A(I14857), .ZN(g6911) );
INV_X32 U_I14860 ( .A(g626), .ZN(I14860) );
INV_X32 U_g6912 ( .A(I14860), .ZN(g6912) );
INV_X32 U_g6942 ( .A(g279), .ZN(g6942) );
INV_X32 U_g6943 ( .A(g801), .ZN(g6943) );
INV_X32 U_I14865 ( .A(g1237), .ZN(I14865) );
INV_X32 U_g6944 ( .A(I14865), .ZN(g6944) );
INV_X32 U_I14868 ( .A(g1237), .ZN(I14868) );
INV_X32 U_g6945 ( .A(I14868), .ZN(g6945) );
INV_X32 U_g6974 ( .A(g1151), .ZN(g6974) );
INV_X32 U_g6977 ( .A(g1145), .ZN(g6977) );
INV_X32 U_g6978 ( .A(g1245), .ZN(g6978) );
INV_X32 U_I14874 ( .A(g1309), .ZN(I14874) );
INV_X32 U_g6979 ( .A(I14874), .ZN(g6979) );
INV_X32 U_I14877 ( .A(g1309), .ZN(I14877) );
INV_X32 U_g6980 ( .A(I14877), .ZN(g6980) );
INV_X32 U_g7009 ( .A(g1352), .ZN(g7009) );
INV_X32 U_g7013 ( .A(g968), .ZN(g7013) );
INV_X32 U_I14882 ( .A(g1786), .ZN(I14882) );
INV_X32 U_g7014 ( .A(I14882), .ZN(g7014) );
INV_X32 U_I14885 ( .A(g1786), .ZN(I14885) );
INV_X32 U_g7015 ( .A(I14885), .ZN(g7015) );
INV_X32 U_I14888 ( .A(g1925), .ZN(I14888) );
INV_X32 U_g7052 ( .A(I14888), .ZN(g7052) );
INV_X32 U_I14891 ( .A(g1925), .ZN(I14891) );
INV_X32 U_g7053 ( .A(I14891), .ZN(g7053) );
INV_X32 U_g7078 ( .A(g1924), .ZN(g7078) );
INV_X32 U_g7079 ( .A(g2040), .ZN(g7079) );
INV_X32 U_g7083 ( .A(g1664), .ZN(g7083) );
INV_X32 U_I14897 ( .A(g2211), .ZN(I14897) );
INV_X32 U_g7084 ( .A(I14897), .ZN(g7084) );
INV_X32 U_I14900 ( .A(g2211), .ZN(I14900) );
INV_X32 U_g7085 ( .A(I14900), .ZN(g7085) );
INV_X32 U_g7134 ( .A(g2727), .ZN(g7134) );
INV_X32 U_g7138 ( .A(g2360), .ZN(g7138) );
INV_X32 U_g7139 ( .A(g1481), .ZN(g7139) );
INV_X32 U_g7140 ( .A(g2170), .ZN(g7140) );
INV_X32 U_g7141 ( .A(g2195), .ZN(g7141) );
INV_X32 U_g7142 ( .A(g8), .ZN(g7142) );
INV_X32 U_g7143 ( .A(g2998), .ZN(g7143) );
INV_X32 U_g7146 ( .A(g3013), .ZN(g7146) );
INV_X32 U_g7149 ( .A(g3105), .ZN(g7149) );
INV_X32 U_g7152 ( .A(g3136), .ZN(g7152) );
INV_X32 U_g7153 ( .A(g480), .ZN(g7153) );
INV_X32 U_g7156 ( .A(g461), .ZN(g7156) );
INV_X32 U_g7157 ( .A(g453), .ZN(g7157) );
INV_X32 U_g7158 ( .A(g1171), .ZN(g7158) );
INV_X32 U_I14917 ( .A(g1312), .ZN(I14917) );
INV_X32 U_g7161 ( .A(I14917), .ZN(g7161) );
INV_X32 U_I14920 ( .A(g1312), .ZN(I14920) );
INV_X32 U_g7162 ( .A(I14920), .ZN(g7162) );
INV_X32 U_g7192 ( .A(g966), .ZN(g7192) );
INV_X32 U_g7193 ( .A(g1491), .ZN(g7193) );
INV_X32 U_I14925 ( .A(g1931), .ZN(I14925) );
INV_X32 U_g7194 ( .A(I14925), .ZN(g7194) );
INV_X32 U_I14928 ( .A(g1931), .ZN(I14928) );
INV_X32 U_g7195 ( .A(I14928), .ZN(g7195) );
INV_X32 U_g7224 ( .A(g1845), .ZN(g7224) );
INV_X32 U_g7227 ( .A(g1839), .ZN(g7227) );
INV_X32 U_g7228 ( .A(g1939), .ZN(g7228) );
INV_X32 U_I14934 ( .A(g2003), .ZN(I14934) );
INV_X32 U_g7229 ( .A(I14934), .ZN(g7229) );
INV_X32 U_I14937 ( .A(g2003), .ZN(I14937) );
INV_X32 U_g7230 ( .A(I14937), .ZN(g7230) );
INV_X32 U_g7259 ( .A(g2046), .ZN(g7259) );
INV_X32 U_g7263 ( .A(g1662), .ZN(g7263) );
INV_X32 U_I14942 ( .A(g2480), .ZN(I14942) );
INV_X32 U_g7264 ( .A(I14942), .ZN(g7264) );
INV_X32 U_I14945 ( .A(g2480), .ZN(I14945) );
INV_X32 U_g7265 ( .A(I14945), .ZN(g7265) );
INV_X32 U_I14948 ( .A(g2619), .ZN(I14948) );
INV_X32 U_g7302 ( .A(I14948), .ZN(g7302) );
INV_X32 U_I14951 ( .A(g2619), .ZN(I14951) );
INV_X32 U_g7303 ( .A(I14951), .ZN(g7303) );
INV_X32 U_g7328 ( .A(g2618), .ZN(g7328) );
INV_X32 U_g7329 ( .A(g2734), .ZN(g7329) );
INV_X32 U_g7333 ( .A(g2358), .ZN(g7333) );
INV_X32 U_I14957 ( .A(g2827), .ZN(I14957) );
INV_X32 U_g7334 ( .A(I14957), .ZN(g7334) );
INV_X32 U_g7335 ( .A(g2827), .ZN(g7335) );
INV_X32 U_g7336 ( .A(g1476), .ZN(g7336) );
INV_X32 U_g7337 ( .A(g2190), .ZN(g7337) );
INV_X32 U_g7338 ( .A(g3002), .ZN(g7338) );
INV_X32 U_g7342 ( .A(g3024), .ZN(g7342) );
INV_X32 U_g7345 ( .A(g3139), .ZN(g7345) );
INV_X32 U_g7346 ( .A(g97), .ZN(g7346) );
INV_X32 U_g7347 ( .A(g490), .ZN(g7347) );
INV_X32 U_g7348 ( .A(g451), .ZN(g7348) );
INV_X32 U_g7349 ( .A(g1167), .ZN(g7349) );
INV_X32 U_g7352 ( .A(g1148), .ZN(g7352) );
INV_X32 U_g7353 ( .A(g1140), .ZN(g7353) );
INV_X32 U_g7354 ( .A(g1865), .ZN(g7354) );
INV_X32 U_I14973 ( .A(g2006), .ZN(I14973) );
INV_X32 U_g7357 ( .A(I14973), .ZN(g7357) );
INV_X32 U_I14976 ( .A(g2006), .ZN(I14976) );
INV_X32 U_g7358 ( .A(I14976), .ZN(g7358) );
INV_X32 U_g7388 ( .A(g1660), .ZN(g7388) );
INV_X32 U_g7389 ( .A(g2185), .ZN(g7389) );
INV_X32 U_I14981 ( .A(g2625), .ZN(I14981) );
INV_X32 U_g7390 ( .A(I14981), .ZN(g7390) );
INV_X32 U_I14984 ( .A(g2625), .ZN(I14984) );
INV_X32 U_g7391 ( .A(I14984), .ZN(g7391) );
INV_X32 U_g7420 ( .A(g2539), .ZN(g7420) );
INV_X32 U_g7423 ( .A(g2533), .ZN(g7423) );
INV_X32 U_g7424 ( .A(g2633), .ZN(g7424) );
INV_X32 U_I14990 ( .A(g2697), .ZN(I14990) );
INV_X32 U_g7425 ( .A(I14990), .ZN(g7425) );
INV_X32 U_I14993 ( .A(g2697), .ZN(I14993) );
INV_X32 U_g7426 ( .A(I14993), .ZN(g7426) );
INV_X32 U_g7455 ( .A(g2740), .ZN(g7455) );
INV_X32 U_g7459 ( .A(g2356), .ZN(g7459) );
INV_X32 U_g7460 ( .A(g1471), .ZN(g7460) );
INV_X32 U_g7461 ( .A(g2175), .ZN(g7461) );
INV_X32 U_g7462 ( .A(g2912), .ZN(g7462) );
INV_X32 U_g7465 ( .A(g2), .ZN(g7465) );
INV_X32 U_g7466 ( .A(g3010), .ZN(g7466) );
INV_X32 U_g7471 ( .A(g3036), .ZN(g7471) );
INV_X32 U_g7475 ( .A(g493), .ZN(g7475) );
INV_X32 U_g7476 ( .A(g785), .ZN(g7476) );
INV_X32 U_g7477 ( .A(g1177), .ZN(g7477) );
INV_X32 U_g7478 ( .A(g1138), .ZN(g7478) );
INV_X32 U_g7479 ( .A(g1861), .ZN(g7479) );
INV_X32 U_g7482 ( .A(g1842), .ZN(g7482) );
INV_X32 U_g7483 ( .A(g1834), .ZN(g7483) );
INV_X32 U_g7484 ( .A(g2559), .ZN(g7484) );
INV_X32 U_I15012 ( .A(g2700), .ZN(I15012) );
INV_X32 U_g7487 ( .A(I15012), .ZN(g7487) );
INV_X32 U_I15015 ( .A(g2700), .ZN(I15015) );
INV_X32 U_g7488 ( .A(I15015), .ZN(g7488) );
INV_X32 U_g7518 ( .A(g2354), .ZN(g7518) );
INV_X32 U_I15019 ( .A(g2830), .ZN(I15019) );
INV_X32 U_g7519 ( .A(I15019), .ZN(g7519) );
INV_X32 U_g7520 ( .A(g2830), .ZN(g7520) );
INV_X32 U_g7521 ( .A(g2200), .ZN(g7521) );
INV_X32 U_g7522 ( .A(g2917), .ZN(g7522) );
INV_X32 U_g7527 ( .A(g3018), .ZN(g7527) );
INV_X32 U_g7529 ( .A(g465), .ZN(g7529) );
INV_X32 U_g7530 ( .A(g496), .ZN(g7530) );
INV_X32 U_g7531 ( .A(g1180), .ZN(g7531) );
INV_X32 U_g7532 ( .A(g1471), .ZN(g7532) );
INV_X32 U_g7533 ( .A(g1871), .ZN(g7533) );
INV_X32 U_g7534 ( .A(g1832), .ZN(g7534) );
INV_X32 U_g7535 ( .A(g2555), .ZN(g7535) );
INV_X32 U_g7538 ( .A(g2536), .ZN(g7538) );
INV_X32 U_g7539 ( .A(g2528), .ZN(g7539) );
INV_X32 U_g7540 ( .A(g1506), .ZN(g7540) );
INV_X32 U_g7541 ( .A(g2180), .ZN(g7541) );
INV_X32 U_g7542 ( .A(g2883), .ZN(g7542) );
INV_X32 U_g7545 ( .A(g2920), .ZN(g7545) );
INV_X32 U_g7548 ( .A(g2990), .ZN(g7548) );
INV_X32 U_g7549 ( .A(g3028), .ZN(g7549) );
INV_X32 U_g7553 ( .A(g3114), .ZN(g7553) );
INV_X32 U_g7554 ( .A(g117), .ZN(g7554) );
INV_X32 U_g7555 ( .A(g1152), .ZN(g7555) );
INV_X32 U_g7556 ( .A(g1183), .ZN(g7556) );
INV_X32 U_g7557 ( .A(g1874), .ZN(g7557) );
INV_X32 U_g7558 ( .A(g2165), .ZN(g7558) );
INV_X32 U_g7559 ( .A(g2565), .ZN(g7559) );
INV_X32 U_g7560 ( .A(g2526), .ZN(g7560) );
INV_X32 U_g7561 ( .A(g1501), .ZN(g7561) );
INV_X32 U_g7562 ( .A(g2888), .ZN(g7562) );
INV_X32 U_g7566 ( .A(g2896), .ZN(g7566) );
INV_X32 U_g7570 ( .A(g3032), .ZN(g7570) );
INV_X32 U_g7573 ( .A(g3120), .ZN(g7573) );
INV_X32 U_g7574 ( .A(g3128), .ZN(g7574) );
INV_X32 U_g7576 ( .A(g468), .ZN(g7576) );
INV_X32 U_g7577 ( .A(g805), .ZN(g7577) );
INV_X32 U_g7578 ( .A(g1846), .ZN(g7578) );
INV_X32 U_g7579 ( .A(g1877), .ZN(g7579) );
INV_X32 U_g7580 ( .A(g2568), .ZN(g7580) );
INV_X32 U_g7581 ( .A(g1496), .ZN(g7581) );
INV_X32 U_g7582 ( .A(g2185), .ZN(g7582) );
INV_X32 U_g7583 ( .A(g2892), .ZN(g7583) );
INV_X32 U_g7587 ( .A(g2903), .ZN(g7587) );
INV_X32 U_g7590 ( .A(g1155), .ZN(g7590) );
INV_X32 U_g7591 ( .A(g1496), .ZN(g7591) );
INV_X32 U_g7592 ( .A(g2540), .ZN(g7592) );
INV_X32 U_g7593 ( .A(g2571), .ZN(g7593) );
INV_X32 U_g7594 ( .A(g2165), .ZN(g7594) );
INV_X32 U_g7595 ( .A(g2900), .ZN(g7595) );
INV_X32 U_g7600 ( .A(g2908), .ZN(g7600) );
INV_X32 U_g7603 ( .A(g3133), .ZN(g7603) );
INV_X32 U_g7604 ( .A(g471), .ZN(g7604) );
INV_X32 U_g7605 ( .A(g1849), .ZN(g7605) );
INV_X32 U_g7606 ( .A(g2190), .ZN(g7606) );
INV_X32 U_g7607 ( .A(g2924), .ZN(g7607) );
INV_X32 U_g7610 ( .A(g312), .ZN(g7610) );
INV_X32 U_g7613 ( .A(g1158), .ZN(g7613) );
INV_X32 U_g7614 ( .A(g2543), .ZN(g7614) );
INV_X32 U_g7615 ( .A(g3123), .ZN(g7615) );
INV_X32 U_g7616 ( .A(g313), .ZN(g7616) );
INV_X32 U_g7619 ( .A(g999), .ZN(g7619) );
INV_X32 U_g7622 ( .A(g1852), .ZN(g7622) );
INV_X32 U_g7623 ( .A(g314), .ZN(g7623) );
INV_X32 U_g7626 ( .A(g315), .ZN(g7626) );
INV_X32 U_g7629 ( .A(g403), .ZN(g7629) );
INV_X32 U_g7632 ( .A(g1000), .ZN(g7632) );
INV_X32 U_g7635 ( .A(g1693), .ZN(g7635) );
INV_X32 U_g7638 ( .A(g2546), .ZN(g7638) );
INV_X32 U_g7639 ( .A(g3094), .ZN(g7639) );
INV_X32 U_g7642 ( .A(g3125), .ZN(g7642) );
INV_X32 U_g7643 ( .A(g316), .ZN(g7643) );
INV_X32 U_g7646 ( .A(g318), .ZN(g7646) );
INV_X32 U_g7649 ( .A(g404), .ZN(g7649) );
INV_X32 U_g7652 ( .A(g1001), .ZN(g7652) );
INV_X32 U_g7655 ( .A(g1002), .ZN(g7655) );
INV_X32 U_g7658 ( .A(g1090), .ZN(g7658) );
INV_X32 U_g7661 ( .A(g1694), .ZN(g7661) );
INV_X32 U_g7664 ( .A(g2387), .ZN(g7664) );
INV_X32 U_g7667 ( .A(g3095), .ZN(g7667) );
INV_X32 U_g7670 ( .A(g317), .ZN(g7670) );
INV_X32 U_g7673 ( .A(g319), .ZN(g7673) );
INV_X32 U_g7676 ( .A(g402), .ZN(g7676) );
INV_X32 U_g7679 ( .A(g1003), .ZN(g7679) );
INV_X32 U_g7682 ( .A(g1005), .ZN(g7682) );
INV_X32 U_g7685 ( .A(g1091), .ZN(g7685) );
INV_X32 U_g7688 ( .A(g1695), .ZN(g7688) );
INV_X32 U_g7691 ( .A(g1696), .ZN(g7691) );
INV_X32 U_g7694 ( .A(g1784), .ZN(g7694) );
INV_X32 U_g7697 ( .A(g2388), .ZN(g7697) );
INV_X32 U_g7700 ( .A(g3096), .ZN(g7700) );
INV_X32 U_g7703 ( .A(g320), .ZN(g7703) );
INV_X32 U_g7706 ( .A(g1004), .ZN(g7706) );
INV_X32 U_g7709 ( .A(g1006), .ZN(g7709) );
INV_X32 U_g7712 ( .A(g1089), .ZN(g7712) );
INV_X32 U_g7715 ( .A(g1697), .ZN(g7715) );
INV_X32 U_g7718 ( .A(g1699), .ZN(g7718) );
INV_X32 U_g7721 ( .A(g1785), .ZN(g7721) );
INV_X32 U_g7724 ( .A(g2389), .ZN(g7724) );
INV_X32 U_g7727 ( .A(g2390), .ZN(g7727) );
INV_X32 U_g7730 ( .A(g2478), .ZN(g7730) );
INV_X32 U_g7733 ( .A(g1007), .ZN(g7733) );
INV_X32 U_g7736 ( .A(g1698), .ZN(g7736) );
INV_X32 U_g7739 ( .A(g1700), .ZN(g7739) );
INV_X32 U_g7742 ( .A(g1783), .ZN(g7742) );
INV_X32 U_g7745 ( .A(g2391), .ZN(g7745) );
INV_X32 U_g7748 ( .A(g2393), .ZN(g7748) );
INV_X32 U_g7751 ( .A(g2479), .ZN(g7751) );
INV_X32 U_g7754 ( .A(g322), .ZN(g7754) );
INV_X32 U_g7757 ( .A(g1701), .ZN(g7757) );
INV_X32 U_g7760 ( .A(g2392), .ZN(g7760) );
INV_X32 U_g7763 ( .A(g2394), .ZN(g7763) );
INV_X32 U_g7766 ( .A(g2477), .ZN(g7766) );
INV_X32 U_g7769 ( .A(g323), .ZN(g7769) );
INV_X32 U_g7772 ( .A(g659), .ZN(g7772) );
INV_X32 U_g7776 ( .A(g1009), .ZN(g7776) );
INV_X32 U_g7779 ( .A(g2395), .ZN(g7779) );
INV_X32 U_g7782 ( .A(g321), .ZN(g7782) );
INV_X32 U_g7785 ( .A(g1010), .ZN(g7785) );
INV_X32 U_g7788 ( .A(g1345), .ZN(g7788) );
INV_X32 U_g7792 ( .A(g1703), .ZN(g7792) );
INV_X32 U_g7796 ( .A(g1008), .ZN(g7796) );
INV_X32 U_g7799 ( .A(g1704), .ZN(g7799) );
INV_X32 U_g7802 ( .A(g2039), .ZN(g7802) );
INV_X32 U_g7806 ( .A(g2397), .ZN(g7806) );
INV_X32 U_g7809 ( .A(g1702), .ZN(g7809) );
INV_X32 U_g7812 ( .A(g2398), .ZN(g7812) );
INV_X32 U_g7815 ( .A(g2733), .ZN(g7815) );
INV_X32 U_g7819 ( .A(g479), .ZN(g7819) );
INV_X32 U_g7822 ( .A(g510), .ZN(g7822) );
INV_X32 U_g7823 ( .A(g2396), .ZN(g7823) );
INV_X32 U_g7826 ( .A(g2987), .ZN(g7826) );
INV_X32 U_g7827 ( .A(g478), .ZN(g7827) );
INV_X32 U_g7830 ( .A(g1166), .ZN(g7830) );
INV_X32 U_g7833 ( .A(g1196), .ZN(g7833) );
INV_X32 U_g7834 ( .A(g2953), .ZN(g7834) );
INV_X32 U_g7837 ( .A(g3044), .ZN(g7837) );
INV_X32 U_g7838 ( .A(g477), .ZN(g7838) );
INV_X32 U_g7841 ( .A(g630), .ZN(g7841) );
INV_X32 U_g7842 ( .A(g1165), .ZN(g7842) );
INV_X32 U_g7845 ( .A(g1860), .ZN(g7845) );
INV_X32 U_g7848 ( .A(g1890), .ZN(g7848) );
INV_X32 U_g7849 ( .A(g2956), .ZN(g7849) );
INV_X32 U_g7852 ( .A(g2981), .ZN(g7852) );
INV_X32 U_g7856 ( .A(g3045), .ZN(g7856) );
INV_X32 U_g7857 ( .A(g3055), .ZN(g7857) );
INV_X32 U_g7858 ( .A(g1164), .ZN(g7858) );
INV_X32 U_g7861 ( .A(g1316), .ZN(g7861) );
INV_X32 U_g7862 ( .A(g1859), .ZN(g7862) );
INV_X32 U_g7865 ( .A(g2554), .ZN(g7865) );
INV_X32 U_g7868 ( .A(g2584), .ZN(g7868) );
INV_X32 U_g7869 ( .A(g2959), .ZN(g7869) );
INV_X32 U_g7872 ( .A(g2874), .ZN(g7872) );
INV_X32 U_g7877 ( .A(g3046), .ZN(g7877) );
INV_X32 U_g7878 ( .A(g3056), .ZN(g7878) );
INV_X32 U_g7879 ( .A(g3065), .ZN(g7879) );
INV_X32 U_g7880 ( .A(g3201), .ZN(g7880) );
INV_X32 U_g7888 ( .A(g1858), .ZN(g7888) );
INV_X32 U_g7891 ( .A(g2010), .ZN(g7891) );
INV_X32 U_g7892 ( .A(g2553), .ZN(g7892) );
INV_X32 U_g7897 ( .A(g3047), .ZN(g7897) );
INV_X32 U_g7898 ( .A(g3057), .ZN(g7898) );
INV_X32 U_g7899 ( .A(g3066), .ZN(g7899) );
INV_X32 U_g7900 ( .A(g3075), .ZN(g7900) );
INV_X32 U_I15222 ( .A(g3151), .ZN(I15222) );
INV_X32 U_g7901 ( .A(I15222), .ZN(g7901) );
INV_X32 U_g7906 ( .A(g488), .ZN(g7906) );
INV_X32 U_I15226 ( .A(g474), .ZN(I15226) );
INV_X32 U_g7909 ( .A(I15226), .ZN(g7909) );
INV_X32 U_g7910 ( .A(g474), .ZN(g7910) );
INV_X32 U_I15230 ( .A(g499), .ZN(I15230) );
INV_X32 U_g7911 ( .A(I15230), .ZN(g7911) );
INV_X32 U_g7912 ( .A(g2552), .ZN(g7912) );
INV_X32 U_g7915 ( .A(g2704), .ZN(g7915) );
INV_X32 U_g7916 ( .A(g2935), .ZN(g7916) );
INV_X32 U_g7919 ( .A(g2963), .ZN(g7919) );
INV_X32 U_g7924 ( .A(g3048), .ZN(g7924) );
INV_X32 U_g7925 ( .A(g3058), .ZN(g7925) );
INV_X32 U_g7926 ( .A(g3067), .ZN(g7926) );
INV_X32 U_g7927 ( .A(g3076), .ZN(g7927) );
INV_X32 U_g7928 ( .A(g3204), .ZN(g7928) );
INV_X32 U_I15256 ( .A(g2950), .ZN(I15256) );
INV_X32 U_g7936 ( .A(I15256), .ZN(g7936) );
INV_X32 U_g7949 ( .A(g165), .ZN(g7949) );
INV_X32 U_g7950 ( .A(g142), .ZN(g7950) );
INV_X32 U_g7953 ( .A(g487), .ZN(g7953) );
INV_X32 U_I15262 ( .A(g481), .ZN(I15262) );
INV_X32 U_g7956 ( .A(I15262), .ZN(g7956) );
INV_X32 U_g7957 ( .A(g481), .ZN(g7957) );
INV_X32 U_g7958 ( .A(g1175), .ZN(g7958) );
INV_X32 U_I15267 ( .A(g1161), .ZN(I15267) );
INV_X32 U_g7961 ( .A(I15267), .ZN(g7961) );
INV_X32 U_g7962 ( .A(g1161), .ZN(g7962) );
INV_X32 U_I15271 ( .A(g1186), .ZN(I15271) );
INV_X32 U_g7963 ( .A(I15271), .ZN(g7963) );
INV_X32 U_g7964 ( .A(g2938), .ZN(g7964) );
INV_X32 U_g7967 ( .A(g2966), .ZN(g7967) );
INV_X32 U_g7971 ( .A(g3049), .ZN(g7971) );
INV_X32 U_g7972 ( .A(g3059), .ZN(g7972) );
INV_X32 U_g7973 ( .A(g3068), .ZN(g7973) );
INV_X32 U_g7974 ( .A(g3077), .ZN(g7974) );
INV_X32 U_g7975 ( .A(g39), .ZN(g7975) );
INV_X32 U_I15288 ( .A(g3109), .ZN(I15288) );
INV_X32 U_g7976 ( .A(I15288), .ZN(g7976) );
INV_X32 U_g7989 ( .A(g3191), .ZN(g7989) );
INV_X32 U_g7990 ( .A(g143), .ZN(g7990) );
INV_X32 U_g7993 ( .A(g145), .ZN(g7993) );
INV_X32 U_g7996 ( .A(g486), .ZN(g7996) );
INV_X32 U_g7999 ( .A(g485), .ZN(g7999) );
INV_X32 U_g8000 ( .A(g853), .ZN(g8000) );
INV_X32 U_g8001 ( .A(g830), .ZN(g8001) );
INV_X32 U_g8004 ( .A(g1174), .ZN(g8004) );
INV_X32 U_I15299 ( .A(g1168), .ZN(I15299) );
INV_X32 U_g8007 ( .A(I15299), .ZN(g8007) );
INV_X32 U_g8008 ( .A(g1168), .ZN(g8008) );
INV_X32 U_g8009 ( .A(g1869), .ZN(g8009) );
INV_X32 U_I15304 ( .A(g1855), .ZN(I15304) );
INV_X32 U_g8012 ( .A(I15304), .ZN(g8012) );
INV_X32 U_g8013 ( .A(g1855), .ZN(g8013) );
INV_X32 U_I15308 ( .A(g1880), .ZN(I15308) );
INV_X32 U_g8014 ( .A(I15308), .ZN(g8014) );
INV_X32 U_g8015 ( .A(g2941), .ZN(g8015) );
INV_X32 U_g8018 ( .A(g2969), .ZN(g8018) );
INV_X32 U_I15313 ( .A(g2930), .ZN(I15313) );
INV_X32 U_g8021 ( .A(I15313), .ZN(g8021) );
INV_X32 U_g8022 ( .A(g2930), .ZN(g8022) );
INV_X32 U_I15317 ( .A(g2842), .ZN(I15317) );
INV_X32 U_g8023 ( .A(I15317), .ZN(g8023) );
INV_X32 U_g8024 ( .A(g2842), .ZN(g8024) );
INV_X32 U_g8025 ( .A(g3050), .ZN(g8025) );
INV_X32 U_g8026 ( .A(g3060), .ZN(g8026) );
INV_X32 U_g8027 ( .A(g3069), .ZN(g8027) );
INV_X32 U_g8028 ( .A(g3078), .ZN(g8028) );
INV_X32 U_g8029 ( .A(g3083), .ZN(g8029) );
INV_X32 U_I15326 ( .A(g3117), .ZN(I15326) );
INV_X32 U_g8030 ( .A(I15326), .ZN(g8030) );
INV_X32 U_I15329 ( .A(g3117), .ZN(I15329) );
INV_X32 U_g8031 ( .A(I15329), .ZN(g8031) );
INV_X32 U_g8044 ( .A(g3194), .ZN(g8044) );
INV_X32 U_g8045 ( .A(g3207), .ZN(g8045) );
INV_X32 U_g8053 ( .A(g141), .ZN(g8053) );
INV_X32 U_g8056 ( .A(g146), .ZN(g8056) );
INV_X32 U_g8059 ( .A(g148), .ZN(g8059) );
INV_X32 U_g8062 ( .A(g169), .ZN(g8062) );
INV_X32 U_g8065 ( .A(g831), .ZN(g8065) );
INV_X32 U_g8068 ( .A(g833), .ZN(g8068) );
INV_X32 U_g8071 ( .A(g1173), .ZN(g8071) );
INV_X32 U_g8074 ( .A(g1172), .ZN(g8074) );
INV_X32 U_g8075 ( .A(g1547), .ZN(g8075) );
INV_X32 U_g8076 ( .A(g1524), .ZN(g8076) );
INV_X32 U_g8079 ( .A(g1868), .ZN(g8079) );
INV_X32 U_I15345 ( .A(g1862), .ZN(I15345) );
INV_X32 U_g8082 ( .A(I15345), .ZN(g8082) );
INV_X32 U_g8083 ( .A(g1862), .ZN(g8083) );
INV_X32 U_g8084 ( .A(g2563), .ZN(g8084) );
INV_X32 U_I15350 ( .A(g2549), .ZN(I15350) );
INV_X32 U_g8087 ( .A(I15350), .ZN(g8087) );
INV_X32 U_g8088 ( .A(g2549), .ZN(g8088) );
INV_X32 U_I15354 ( .A(g2574), .ZN(I15354) );
INV_X32 U_g8089 ( .A(I15354), .ZN(g8089) );
INV_X32 U_g8090 ( .A(g2944), .ZN(g8090) );
INV_X32 U_g8093 ( .A(g2972), .ZN(g8093) );
INV_X32 U_I15359 ( .A(g2858), .ZN(I15359) );
INV_X32 U_g8096 ( .A(I15359), .ZN(g8096) );
INV_X32 U_g8097 ( .A(g2858), .ZN(g8097) );
INV_X32 U_g8098 ( .A(g3051), .ZN(g8098) );
INV_X32 U_g8099 ( .A(g3061), .ZN(g8099) );
INV_X32 U_g8100 ( .A(g3070), .ZN(g8100) );
INV_X32 U_g8101 ( .A(g2997), .ZN(g8101) );
INV_X32 U_g8102 ( .A(g27), .ZN(g8102) );
INV_X32 U_g8103 ( .A(g185), .ZN(g8103) );
INV_X32 U_I15369 ( .A(g3129), .ZN(I15369) );
INV_X32 U_g8106 ( .A(I15369), .ZN(g8106) );
INV_X32 U_I15372 ( .A(g3129), .ZN(I15372) );
INV_X32 U_g8107 ( .A(I15372), .ZN(g8107) );
INV_X32 U_g8120 ( .A(g3197), .ZN(g8120) );
INV_X32 U_g8123 ( .A(g144), .ZN(g8123) );
INV_X32 U_g8126 ( .A(g149), .ZN(g8126) );
INV_X32 U_g8129 ( .A(g151), .ZN(g8129) );
INV_X32 U_g8132 ( .A(g170), .ZN(g8132) );
INV_X32 U_g8135 ( .A(g172), .ZN(g8135) );
INV_X32 U_g8138 ( .A(g829), .ZN(g8138) );
INV_X32 U_g8141 ( .A(g834), .ZN(g8141) );
INV_X32 U_g8144 ( .A(g836), .ZN(g8144) );
INV_X32 U_g8147 ( .A(g857), .ZN(g8147) );
INV_X32 U_g8150 ( .A(g1525), .ZN(g8150) );
INV_X32 U_g8153 ( .A(g1527), .ZN(g8153) );
INV_X32 U_g8156 ( .A(g1867), .ZN(g8156) );
INV_X32 U_g8159 ( .A(g1866), .ZN(g8159) );
INV_X32 U_g8160 ( .A(g2241), .ZN(g8160) );
INV_X32 U_g8161 ( .A(g2218), .ZN(g8161) );
INV_X32 U_g8164 ( .A(g2562), .ZN(g8164) );
INV_X32 U_I15392 ( .A(g2556), .ZN(I15392) );
INV_X32 U_g8167 ( .A(I15392), .ZN(g8167) );
INV_X32 U_g8168 ( .A(g2556), .ZN(g8168) );
INV_X32 U_g8169 ( .A(g2947), .ZN(g8169) );
INV_X32 U_g8172 ( .A(g2975), .ZN(g8172) );
INV_X32 U_I15398 ( .A(g2845), .ZN(I15398) );
INV_X32 U_g8175 ( .A(I15398), .ZN(g8175) );
INV_X32 U_g8176 ( .A(g2845), .ZN(g8176) );
INV_X32 U_g8177 ( .A(g3043), .ZN(g8177) );
INV_X32 U_g8178 ( .A(g3052), .ZN(g8178) );
INV_X32 U_g8179 ( .A(g3062), .ZN(g8179) );
INV_X32 U_g8180 ( .A(g3071), .ZN(g8180) );
INV_X32 U_g8181 ( .A(g48), .ZN(g8181) );
INV_X32 U_g8182 ( .A(g3198), .ZN(g8182) );
INV_X32 U_g8183 ( .A(g3188), .ZN(g8183) );
INV_X32 U_g8191 ( .A(g147), .ZN(g8191) );
INV_X32 U_g8194 ( .A(g152), .ZN(g8194) );
INV_X32 U_g8197 ( .A(g154), .ZN(g8197) );
INV_X32 U_g8200 ( .A(g168), .ZN(g8200) );
INV_X32 U_g8203 ( .A(g173), .ZN(g8203) );
INV_X32 U_g8206 ( .A(g175), .ZN(g8206) );
INV_X32 U_g8209 ( .A(g832), .ZN(g8209) );
INV_X32 U_g8212 ( .A(g837), .ZN(g8212) );
INV_X32 U_g8215 ( .A(g839), .ZN(g8215) );
INV_X32 U_g8218 ( .A(g858), .ZN(g8218) );
INV_X32 U_g8221 ( .A(g860), .ZN(g8221) );
INV_X32 U_g8224 ( .A(g1523), .ZN(g8224) );
INV_X32 U_g8227 ( .A(g1528), .ZN(g8227) );
INV_X32 U_g8230 ( .A(g1530), .ZN(g8230) );
INV_X32 U_g8233 ( .A(g1551), .ZN(g8233) );
INV_X32 U_g8236 ( .A(g2219), .ZN(g8236) );
INV_X32 U_g8239 ( .A(g2221), .ZN(g8239) );
INV_X32 U_g8242 ( .A(g2561), .ZN(g8242) );
INV_X32 U_g8245 ( .A(g2560), .ZN(g8245) );
INV_X32 U_g8246 ( .A(g2978), .ZN(g8246) );
INV_X32 U_I15429 ( .A(g2833), .ZN(I15429) );
INV_X32 U_g8249 ( .A(I15429), .ZN(g8249) );
INV_X32 U_g8250 ( .A(g2833), .ZN(g8250) );
INV_X32 U_I15433 ( .A(g2861), .ZN(I15433) );
INV_X32 U_g8251 ( .A(I15433), .ZN(g8251) );
INV_X32 U_g8252 ( .A(g2861), .ZN(g8252) );
INV_X32 U_g8253 ( .A(g3053), .ZN(g8253) );
INV_X32 U_g8254 ( .A(g3063), .ZN(g8254) );
INV_X32 U_g8255 ( .A(g3072), .ZN(g8255) );
INV_X32 U_g8256 ( .A(g30), .ZN(g8256) );
INV_X32 U_g8257 ( .A(g3201), .ZN(g8257) );
INV_X32 U_I15442 ( .A(g3235), .ZN(I15442) );
INV_X32 U_g8258 ( .A(I15442), .ZN(g8258) );
INV_X32 U_I15445 ( .A(g3236), .ZN(I15445) );
INV_X32 U_g8259 ( .A(I15445), .ZN(g8259) );
INV_X32 U_I15448 ( .A(g3237), .ZN(I15448) );
INV_X32 U_g8260 ( .A(I15448), .ZN(g8260) );
INV_X32 U_I15451 ( .A(g3238), .ZN(I15451) );
INV_X32 U_g8261 ( .A(I15451), .ZN(g8261) );
INV_X32 U_I15454 ( .A(g3239), .ZN(I15454) );
INV_X32 U_g8262 ( .A(I15454), .ZN(g8262) );
INV_X32 U_I15457 ( .A(g3240), .ZN(I15457) );
INV_X32 U_g8263 ( .A(I15457), .ZN(g8263) );
INV_X32 U_I15460 ( .A(g3241), .ZN(I15460) );
INV_X32 U_g8264 ( .A(I15460), .ZN(g8264) );
INV_X32 U_I15463 ( .A(g3242), .ZN(I15463) );
INV_X32 U_g8265 ( .A(I15463), .ZN(g8265) );
INV_X32 U_I15466 ( .A(g3243), .ZN(I15466) );
INV_X32 U_g8266 ( .A(I15466), .ZN(g8266) );
INV_X32 U_I15469 ( .A(g3244), .ZN(I15469) );
INV_X32 U_g8267 ( .A(I15469), .ZN(g8267) );
INV_X32 U_I15472 ( .A(g3245), .ZN(I15472) );
INV_X32 U_g8268 ( .A(I15472), .ZN(g8268) );
INV_X32 U_I15475 ( .A(g3246), .ZN(I15475) );
INV_X32 U_g8269 ( .A(I15475), .ZN(g8269) );
INV_X32 U_I15478 ( .A(g3247), .ZN(I15478) );
INV_X32 U_g8270 ( .A(I15478), .ZN(g8270) );
INV_X32 U_I15481 ( .A(g3248), .ZN(I15481) );
INV_X32 U_g8271 ( .A(I15481), .ZN(g8271) );
INV_X32 U_I15484 ( .A(g3249), .ZN(I15484) );
INV_X32 U_g8272 ( .A(I15484), .ZN(g8272) );
INV_X32 U_I15487 ( .A(g3250), .ZN(I15487) );
INV_X32 U_g8273 ( .A(I15487), .ZN(g8273) );
INV_X32 U_I15490 ( .A(g3251), .ZN(I15490) );
INV_X32 U_g8274 ( .A(I15490), .ZN(g8274) );
INV_X32 U_I15493 ( .A(g3252), .ZN(I15493) );
INV_X32 U_g8275 ( .A(I15493), .ZN(g8275) );
INV_X32 U_g8276 ( .A(g3253), .ZN(g8276) );
INV_X32 U_g8277 ( .A(g3305), .ZN(g8277) );
INV_X32 U_g8278 ( .A(g3337), .ZN(g8278) );
INV_X32 U_I15499 ( .A(g7911), .ZN(I15499) );
INV_X32 U_g8284 ( .A(I15499), .ZN(g8284) );
INV_X32 U_g8285 ( .A(g3365), .ZN(g8285) );
INV_X32 U_g8286 ( .A(g3461), .ZN(g8286) );
INV_X32 U_g8287 ( .A(g3493), .ZN(g8287) );
INV_X32 U_I15505 ( .A(g7963), .ZN(I15505) );
INV_X32 U_g8293 ( .A(I15505), .ZN(g8293) );
INV_X32 U_g8294 ( .A(g3521), .ZN(g8294) );
INV_X32 U_g8295 ( .A(g3617), .ZN(g8295) );
INV_X32 U_g8296 ( .A(g3649), .ZN(g8296) );
INV_X32 U_I15511 ( .A(g8014), .ZN(I15511) );
INV_X32 U_g8302 ( .A(I15511), .ZN(g8302) );
INV_X32 U_g8303 ( .A(g3677), .ZN(g8303) );
INV_X32 U_g8304 ( .A(g3773), .ZN(g8304) );
INV_X32 U_g8305 ( .A(g3805), .ZN(g8305) );
INV_X32 U_I15517 ( .A(g8089), .ZN(I15517) );
INV_X32 U_g8311 ( .A(I15517), .ZN(g8311) );
INV_X32 U_g8312 ( .A(g3833), .ZN(g8312) );
INV_X32 U_g8313 ( .A(g3897), .ZN(g8313) );
INV_X32 U_g8317 ( .A(g3919), .ZN(g8317) );
INV_X32 U_I15523 ( .A(g3254), .ZN(I15523) );
INV_X32 U_g8321 ( .A(I15523), .ZN(g8321) );
INV_X32 U_I15526 ( .A(g6314), .ZN(I15526) );
INV_X32 U_g8324 ( .A(I15526), .ZN(g8324) );
INV_X32 U_I15532 ( .A(g3410), .ZN(I15532) );
INV_X32 U_g8330 ( .A(I15532), .ZN(g8330) );
INV_X32 U_I15535 ( .A(g6519), .ZN(I15535) );
INV_X32 U_g8333 ( .A(I15535), .ZN(g8333) );
INV_X32 U_I15538 ( .A(g6369), .ZN(I15538) );
INV_X32 U_g8336 ( .A(I15538), .ZN(g8336) );
INV_X32 U_I15543 ( .A(g3410), .ZN(I15543) );
INV_X32 U_g8341 ( .A(I15543), .ZN(g8341) );
INV_X32 U_I15546 ( .A(g6783), .ZN(I15546) );
INV_X32 U_g8344 ( .A(I15546), .ZN(g8344) );
INV_X32 U_I15549 ( .A(g6574), .ZN(I15549) );
INV_X32 U_g8347 ( .A(I15549), .ZN(g8347) );
INV_X32 U_I15553 ( .A(g3566), .ZN(I15553) );
INV_X32 U_g8351 ( .A(I15553), .ZN(g8351) );
INV_X32 U_I15556 ( .A(g6783), .ZN(I15556) );
INV_X32 U_g8354 ( .A(I15556), .ZN(g8354) );
INV_X32 U_I15559 ( .A(g7015), .ZN(I15559) );
INV_X32 U_g8357 ( .A(I15559), .ZN(g8357) );
INV_X32 U_I15562 ( .A(g5778), .ZN(I15562) );
INV_X32 U_g8360 ( .A(I15562), .ZN(g8360) );
INV_X32 U_I15565 ( .A(g6838), .ZN(I15565) );
INV_X32 U_g8363 ( .A(I15565), .ZN(g8363) );
INV_X32 U_I15568 ( .A(g3722), .ZN(I15568) );
INV_X32 U_g8366 ( .A(I15568), .ZN(g8366) );
INV_X32 U_I15571 ( .A(g7085), .ZN(I15571) );
INV_X32 U_g8369 ( .A(I15571), .ZN(g8369) );
INV_X32 U_I15574 ( .A(g6838), .ZN(I15574) );
INV_X32 U_g8372 ( .A(I15574), .ZN(g8372) );
INV_X32 U_I15577 ( .A(g7265), .ZN(I15577) );
INV_X32 U_g8375 ( .A(I15577), .ZN(g8375) );
INV_X32 U_I15580 ( .A(g5837), .ZN(I15580) );
INV_X32 U_g8378 ( .A(I15580), .ZN(g8378) );
INV_X32 U_I15584 ( .A(g3254), .ZN(I15584) );
INV_X32 U_g8382 ( .A(I15584), .ZN(g8382) );
INV_X32 U_I15590 ( .A(g3410), .ZN(I15590) );
INV_X32 U_g8388 ( .A(I15590), .ZN(g8388) );
INV_X32 U_I15593 ( .A(g6519), .ZN(I15593) );
INV_X32 U_g8391 ( .A(I15593), .ZN(g8391) );
INV_X32 U_I15599 ( .A(g3566), .ZN(I15599) );
INV_X32 U_g8397 ( .A(I15599), .ZN(g8397) );
INV_X32 U_I15602 ( .A(g6783), .ZN(I15602) );
INV_X32 U_g8400 ( .A(I15602), .ZN(g8400) );
INV_X32 U_I15605 ( .A(g6574), .ZN(I15605) );
INV_X32 U_g8403 ( .A(I15605), .ZN(g8403) );
INV_X32 U_I15610 ( .A(g3566), .ZN(I15610) );
INV_X32 U_g8408 ( .A(I15610), .ZN(g8408) );
INV_X32 U_I15613 ( .A(g7085), .ZN(I15613) );
INV_X32 U_g8411 ( .A(I15613), .ZN(g8411) );
INV_X32 U_I15616 ( .A(g6838), .ZN(I15616) );
INV_X32 U_g8414 ( .A(I15616), .ZN(g8414) );
INV_X32 U_I15620 ( .A(g3722), .ZN(I15620) );
INV_X32 U_g8418 ( .A(I15620), .ZN(g8418) );
INV_X32 U_I15623 ( .A(g7085), .ZN(I15623) );
INV_X32 U_g8421 ( .A(I15623), .ZN(g8421) );
INV_X32 U_I15626 ( .A(g7265), .ZN(I15626) );
INV_X32 U_g8424 ( .A(I15626), .ZN(g8424) );
INV_X32 U_I15629 ( .A(g5837), .ZN(I15629) );
INV_X32 U_g8427 ( .A(I15629), .ZN(g8427) );
INV_X32 U_I15636 ( .A(g3410), .ZN(I15636) );
INV_X32 U_g8434 ( .A(I15636), .ZN(g8434) );
INV_X32 U_I15642 ( .A(g3566), .ZN(I15642) );
INV_X32 U_g8440 ( .A(I15642), .ZN(g8440) );
INV_X32 U_I15645 ( .A(g6783), .ZN(I15645) );
INV_X32 U_g8443 ( .A(I15645), .ZN(g8443) );
INV_X32 U_I15651 ( .A(g3722), .ZN(I15651) );
INV_X32 U_g8449 ( .A(I15651), .ZN(g8449) );
INV_X32 U_I15654 ( .A(g7085), .ZN(I15654) );
INV_X32 U_g8452 ( .A(I15654), .ZN(g8452) );
INV_X32 U_I15657 ( .A(g6838), .ZN(I15657) );
INV_X32 U_g8455 ( .A(I15657), .ZN(g8455) );
INV_X32 U_I15662 ( .A(g3722), .ZN(I15662) );
INV_X32 U_g8460 ( .A(I15662), .ZN(g8460) );
INV_X32 U_I15671 ( .A(g3566), .ZN(I15671) );
INV_X32 U_g8469 ( .A(I15671), .ZN(g8469) );
INV_X32 U_I15677 ( .A(g3722), .ZN(I15677) );
INV_X32 U_g8475 ( .A(I15677), .ZN(g8475) );
INV_X32 U_I15680 ( .A(g7085), .ZN(I15680) );
INV_X32 U_g8478 ( .A(I15680), .ZN(g8478) );
INV_X32 U_I15696 ( .A(g3722), .ZN(I15696) );
INV_X32 U_g8494 ( .A(I15696), .ZN(g8494) );
INV_X32 U_g8514 ( .A(g6139), .ZN(g8514) );
INV_X32 U_g8530 ( .A(g6156), .ZN(g8530) );
INV_X32 U_g8568 ( .A(g6230), .ZN(g8568) );
INV_X32 U_I15771 ( .A(g6000), .ZN(I15771) );
INV_X32 U_g8569 ( .A(I15771), .ZN(g8569) );
INV_X32 U_I15779 ( .A(g6000), .ZN(I15779) );
INV_X32 U_g8575 ( .A(I15779), .ZN(g8575) );
INV_X32 U_I15784 ( .A(g6000), .ZN(I15784) );
INV_X32 U_g8578 ( .A(I15784), .ZN(g8578) );
INV_X32 U_I15787 ( .A(g6000), .ZN(I15787) );
INV_X32 U_g8579 ( .A(I15787), .ZN(g8579) );
INV_X32 U_g8580 ( .A(g6281), .ZN(g8580) );
INV_X32 U_g8587 ( .A(g6418), .ZN(g8587) );
INV_X32 U_g8594 ( .A(g6623), .ZN(g8594) );
INV_X32 U_I15794 ( .A(g3338), .ZN(I15794) );
INV_X32 U_g8602 ( .A(I15794), .ZN(g8602) );
INV_X32 U_g8605 ( .A(g6887), .ZN(g8605) );
INV_X32 U_I15800 ( .A(g3494), .ZN(I15800) );
INV_X32 U_g8614 ( .A(I15800), .ZN(g8614) );
INV_X32 U_I15803 ( .A(g8107), .ZN(I15803) );
INV_X32 U_g8617 ( .A(I15803), .ZN(g8617) );
INV_X32 U_I15806 ( .A(g5550), .ZN(I15806) );
INV_X32 U_g8620 ( .A(I15806), .ZN(g8620) );
INV_X32 U_I15810 ( .A(g3338), .ZN(I15810) );
INV_X32 U_g8622 ( .A(I15810), .ZN(g8622) );
INV_X32 U_I15815 ( .A(g3650), .ZN(I15815) );
INV_X32 U_g8627 ( .A(I15815), .ZN(g8627) );
INV_X32 U_I15818 ( .A(g5596), .ZN(I15818) );
INV_X32 U_g8630 ( .A(I15818), .ZN(g8630) );
INV_X32 U_I15822 ( .A(g3494), .ZN(I15822) );
INV_X32 U_g8632 ( .A(I15822), .ZN(g8632) );
INV_X32 U_I15827 ( .A(g3806), .ZN(I15827) );
INV_X32 U_g8637 ( .A(I15827), .ZN(g8637) );
INV_X32 U_I15830 ( .A(g8031), .ZN(I15830) );
INV_X32 U_g8640 ( .A(I15830), .ZN(g8640) );
INV_X32 U_I15833 ( .A(g3338), .ZN(I15833) );
INV_X32 U_g8643 ( .A(I15833), .ZN(g8643) );
INV_X32 U_I15836 ( .A(g3366), .ZN(I15836) );
INV_X32 U_g8646 ( .A(I15836), .ZN(g8646) );
INV_X32 U_I15839 ( .A(g5613), .ZN(I15839) );
INV_X32 U_g8649 ( .A(I15839), .ZN(g8649) );
INV_X32 U_I15843 ( .A(g3650), .ZN(I15843) );
INV_X32 U_g8651 ( .A(I15843), .ZN(g8651) );
INV_X32 U_I15847 ( .A(g3878), .ZN(I15847) );
INV_X32 U_g8655 ( .A(I15847), .ZN(g8655) );
INV_X32 U_I15850 ( .A(g5627), .ZN(I15850) );
INV_X32 U_g8658 ( .A(I15850), .ZN(g8658) );
INV_X32 U_I15853 ( .A(g3494), .ZN(I15853) );
INV_X32 U_g8659 ( .A(I15853), .ZN(g8659) );
INV_X32 U_I15856 ( .A(g3522), .ZN(I15856) );
INV_X32 U_g8662 ( .A(I15856), .ZN(g8662) );
INV_X32 U_I15859 ( .A(g5638), .ZN(I15859) );
INV_X32 U_g8665 ( .A(I15859), .ZN(g8665) );
INV_X32 U_I15863 ( .A(g3806), .ZN(I15863) );
INV_X32 U_g8667 ( .A(I15863), .ZN(g8667) );
INV_X32 U_I15866 ( .A(g3878), .ZN(I15866) );
INV_X32 U_g8670 ( .A(I15866), .ZN(g8670) );
INV_X32 U_I15869 ( .A(g7976), .ZN(I15869) );
INV_X32 U_g8673 ( .A(I15869), .ZN(g8673) );
INV_X32 U_I15873 ( .A(g5655), .ZN(I15873) );
INV_X32 U_g8677 ( .A(I15873), .ZN(g8677) );
INV_X32 U_I15876 ( .A(g3650), .ZN(I15876) );
INV_X32 U_g8678 ( .A(I15876), .ZN(g8678) );
INV_X32 U_I15879 ( .A(g3678), .ZN(I15879) );
INV_X32 U_g8681 ( .A(I15879), .ZN(g8681) );
INV_X32 U_I15882 ( .A(g3878), .ZN(I15882) );
INV_X32 U_g8684 ( .A(I15882), .ZN(g8684) );
INV_X32 U_I15887 ( .A(g5693), .ZN(I15887) );
INV_X32 U_g8689 ( .A(I15887), .ZN(g8689) );
INV_X32 U_I15890 ( .A(g3806), .ZN(I15890) );
INV_X32 U_g8690 ( .A(I15890), .ZN(g8690) );
INV_X32 U_I15893 ( .A(g3834), .ZN(I15893) );
INV_X32 U_g8693 ( .A(I15893), .ZN(g8693) );
INV_X32 U_I15896 ( .A(g3878), .ZN(I15896) );
INV_X32 U_g8696 ( .A(I15896), .ZN(g8696) );
INV_X32 U_I15899 ( .A(g5626), .ZN(I15899) );
INV_X32 U_g8699 ( .A(I15899), .ZN(g8699) );
INV_X32 U_I15902 ( .A(g6486), .ZN(I15902) );
INV_X32 U_g8700 ( .A(I15902), .ZN(g8700) );
INV_X32 U_I15909 ( .A(g5745), .ZN(I15909) );
INV_X32 U_g8707 ( .A(I15909), .ZN(g8707) );
INV_X32 U_I15912 ( .A(g3878), .ZN(I15912) );
INV_X32 U_g8708 ( .A(I15912), .ZN(g8708) );
INV_X32 U_I15915 ( .A(g3878), .ZN(I15915) );
INV_X32 U_g8711 ( .A(I15915), .ZN(g8711) );
INV_X32 U_I15918 ( .A(g6643), .ZN(I15918) );
INV_X32 U_g8714 ( .A(I15918), .ZN(g8714) );
INV_X32 U_I15922 ( .A(g5654), .ZN(I15922) );
INV_X32 U_g8718 ( .A(I15922), .ZN(g8718) );
INV_X32 U_I15925 ( .A(g6751), .ZN(I15925) );
INV_X32 U_g8719 ( .A(I15925), .ZN(g8719) );
INV_X32 U_I15932 ( .A(g5423), .ZN(I15932) );
INV_X32 U_g8726 ( .A(I15932), .ZN(g8726) );
INV_X32 U_I15935 ( .A(g3878), .ZN(I15935) );
INV_X32 U_g8745 ( .A(I15935), .ZN(g8745) );
INV_X32 U_I15938 ( .A(g3338), .ZN(I15938) );
INV_X32 U_g8748 ( .A(I15938), .ZN(g8748) );
INV_X32 U_I15942 ( .A(g6945), .ZN(I15942) );
INV_X32 U_g8752 ( .A(I15942), .ZN(g8752) );
INV_X32 U_I15946 ( .A(g5692), .ZN(I15946) );
INV_X32 U_g8756 ( .A(I15946), .ZN(g8756) );
INV_X32 U_I15949 ( .A(g7053), .ZN(I15949) );
INV_X32 U_g8757 ( .A(I15949), .ZN(g8757) );
INV_X32 U_I15955 ( .A(g3878), .ZN(I15955) );
INV_X32 U_g8763 ( .A(I15955), .ZN(g8763) );
INV_X32 U_I15958 ( .A(g3878), .ZN(I15958) );
INV_X32 U_g8766 ( .A(I15958), .ZN(g8766) );
INV_X32 U_I15961 ( .A(g6051), .ZN(I15961) );
INV_X32 U_g8769 ( .A(I15961), .ZN(g8769) );
INV_X32 U_I15964 ( .A(g7554), .ZN(I15964) );
INV_X32 U_g8770 ( .A(I15964), .ZN(g8770) );
INV_X32 U_I15967 ( .A(g3494), .ZN(I15967) );
INV_X32 U_g8771 ( .A(I15967), .ZN(g8771) );
INV_X32 U_I15971 ( .A(g7195), .ZN(I15971) );
INV_X32 U_g8775 ( .A(I15971), .ZN(g8775) );
INV_X32 U_I15975 ( .A(g5744), .ZN(I15975) );
INV_X32 U_g8779 ( .A(I15975), .ZN(g8779) );
INV_X32 U_I15978 ( .A(g7303), .ZN(I15978) );
INV_X32 U_g8780 ( .A(I15978), .ZN(g8780) );
INV_X32 U_I15983 ( .A(g3878), .ZN(I15983) );
INV_X32 U_g8785 ( .A(I15983), .ZN(g8785) );
INV_X32 U_I15986 ( .A(g3878), .ZN(I15986) );
INV_X32 U_g8788 ( .A(I15986), .ZN(g8788) );
INV_X32 U_I15989 ( .A(g6053), .ZN(I15989) );
INV_X32 U_g8791 ( .A(I15989), .ZN(g8791) );
INV_X32 U_I15992 ( .A(g6055), .ZN(I15992) );
INV_X32 U_g8792 ( .A(I15992), .ZN(g8792) );
INV_X32 U_I15995 ( .A(g7577), .ZN(I15995) );
INV_X32 U_g8793 ( .A(I15995), .ZN(g8793) );
INV_X32 U_I15998 ( .A(g3650), .ZN(I15998) );
INV_X32 U_g8794 ( .A(I15998), .ZN(g8794) );
INV_X32 U_I16002 ( .A(g7391), .ZN(I16002) );
INV_X32 U_g8798 ( .A(I16002), .ZN(g8798) );
INV_X32 U_I16006 ( .A(g3878), .ZN(I16006) );
INV_X32 U_g8802 ( .A(I16006), .ZN(g8802) );
INV_X32 U_I16009 ( .A(g3878), .ZN(I16009) );
INV_X32 U_g8805 ( .A(I16009), .ZN(g8805) );
INV_X32 U_I16012 ( .A(g5390), .ZN(I16012) );
INV_X32 U_g8808 ( .A(I16012), .ZN(g8808) );
INV_X32 U_I16015 ( .A(g6056), .ZN(I16015) );
INV_X32 U_g8809 ( .A(I16015), .ZN(g8809) );
INV_X32 U_I16018 ( .A(g6058), .ZN(I16018) );
INV_X32 U_g8810 ( .A(I16018), .ZN(g8810) );
INV_X32 U_I16021 ( .A(g6060), .ZN(I16021) );
INV_X32 U_g8811 ( .A(I16021), .ZN(g8811) );
INV_X32 U_I16024 ( .A(g7591), .ZN(I16024) );
INV_X32 U_g8812 ( .A(I16024), .ZN(g8812) );
INV_X32 U_I16027 ( .A(g3806), .ZN(I16027) );
INV_X32 U_g8813 ( .A(I16027), .ZN(g8813) );
INV_X32 U_I16031 ( .A(g3878), .ZN(I16031) );
INV_X32 U_g8817 ( .A(I16031), .ZN(g8817) );
INV_X32 U_I16034 ( .A(g5396), .ZN(I16034) );
INV_X32 U_g8820 ( .A(I16034), .ZN(g8820) );
INV_X32 U_I16037 ( .A(g6061), .ZN(I16037) );
INV_X32 U_g8821 ( .A(I16037), .ZN(g8821) );
INV_X32 U_g8822 ( .A(g4602), .ZN(g8822) );
INV_X32 U_I16041 ( .A(g6486), .ZN(I16041) );
INV_X32 U_g8823 ( .A(I16041), .ZN(g8823) );
INV_X32 U_I16044 ( .A(g5397), .ZN(I16044) );
INV_X32 U_g8824 ( .A(I16044), .ZN(g8824) );
INV_X32 U_I16047 ( .A(g6063), .ZN(I16047) );
INV_X32 U_g8825 ( .A(I16047), .ZN(g8825) );
INV_X32 U_I16050 ( .A(g6065), .ZN(I16050) );
INV_X32 U_g8826 ( .A(I16050), .ZN(g8826) );
INV_X32 U_I16053 ( .A(g6067), .ZN(I16053) );
INV_X32 U_g8827 ( .A(I16053), .ZN(g8827) );
INV_X32 U_I16056 ( .A(g7606), .ZN(I16056) );
INV_X32 U_g8828 ( .A(I16056), .ZN(g8828) );
INV_X32 U_I16059 ( .A(g3878), .ZN(I16059) );
INV_X32 U_g8829 ( .A(I16059), .ZN(g8829) );
INV_X32 U_I16062 ( .A(g3900), .ZN(I16062) );
INV_X32 U_g8832 ( .A(I16062), .ZN(g8832) );
INV_X32 U_I16065 ( .A(g7936), .ZN(I16065) );
INV_X32 U_g8835 ( .A(I16065), .ZN(g8835) );
INV_X32 U_I16068 ( .A(g5438), .ZN(I16068) );
INV_X32 U_g8836 ( .A(I16068), .ZN(g8836) );
INV_X32 U_I16071 ( .A(g5395), .ZN(I16071) );
INV_X32 U_g8839 ( .A(I16071), .ZN(g8839) );
INV_X32 U_I16074 ( .A(g5399), .ZN(I16074) );
INV_X32 U_g8840 ( .A(I16074), .ZN(g8840) );
INV_X32 U_I16079 ( .A(g6086), .ZN(I16079) );
INV_X32 U_g8843 ( .A(I16079), .ZN(g8843) );
INV_X32 U_I16082 ( .A(g5401), .ZN(I16082) );
INV_X32 U_g8844 ( .A(I16082), .ZN(g8844) );
INV_X32 U_I16085 ( .A(g6080), .ZN(I16085) );
INV_X32 U_g8845 ( .A(I16085), .ZN(g8845) );
INV_X32 U_g8846 ( .A(g4779), .ZN(g8846) );
INV_X32 U_I16089 ( .A(g6751), .ZN(I16089) );
INV_X32 U_g8847 ( .A(I16089), .ZN(g8847) );
INV_X32 U_I16092 ( .A(g5402), .ZN(I16092) );
INV_X32 U_g8850 ( .A(I16092), .ZN(g8850) );
INV_X32 U_I16095 ( .A(g6082), .ZN(I16095) );
INV_X32 U_g8851 ( .A(I16095), .ZN(g8851) );
INV_X32 U_I16098 ( .A(g6084), .ZN(I16098) );
INV_X32 U_g8852 ( .A(I16098), .ZN(g8852) );
INV_X32 U_I16101 ( .A(g3878), .ZN(I16101) );
INV_X32 U_g8853 ( .A(I16101), .ZN(g8853) );
INV_X32 U_I16104 ( .A(g6448), .ZN(I16104) );
INV_X32 U_g8856 ( .A(I16104), .ZN(g8856) );
INV_X32 U_I16107 ( .A(g5398), .ZN(I16107) );
INV_X32 U_g8859 ( .A(I16107), .ZN(g8859) );
INV_X32 U_I16110 ( .A(g5404), .ZN(I16110) );
INV_X32 U_g8860 ( .A(I16110), .ZN(g8860) );
INV_X32 U_I16114 ( .A(g7936), .ZN(I16114) );
INV_X32 U_g8862 ( .A(I16114), .ZN(g8862) );
INV_X32 U_I16117 ( .A(g5473), .ZN(I16117) );
INV_X32 U_g8863 ( .A(I16117), .ZN(g8863) );
INV_X32 U_I16120 ( .A(g5400), .ZN(I16120) );
INV_X32 U_g8866 ( .A(I16120), .ZN(g8866) );
INV_X32 U_I16123 ( .A(g5406), .ZN(I16123) );
INV_X32 U_g8867 ( .A(I16123), .ZN(g8867) );
INV_X32 U_I16128 ( .A(g6103), .ZN(I16128) );
INV_X32 U_g8870 ( .A(I16128), .ZN(g8870) );
INV_X32 U_I16131 ( .A(g5408), .ZN(I16131) );
INV_X32 U_g8871 ( .A(I16131), .ZN(g8871) );
INV_X32 U_I16134 ( .A(g6099), .ZN(I16134) );
INV_X32 U_g8872 ( .A(I16134), .ZN(g8872) );
INV_X32 U_g8873 ( .A(g4955), .ZN(g8873) );
INV_X32 U_I16138 ( .A(g7053), .ZN(I16138) );
INV_X32 U_g8874 ( .A(I16138), .ZN(g8874) );
INV_X32 U_I16141 ( .A(g5409), .ZN(I16141) );
INV_X32 U_g8877 ( .A(I16141), .ZN(g8877) );
INV_X32 U_I16144 ( .A(g6101), .ZN(I16144) );
INV_X32 U_g8878 ( .A(I16144), .ZN(g8878) );
INV_X32 U_I16147 ( .A(g3878), .ZN(I16147) );
INV_X32 U_g8879 ( .A(I16147), .ZN(g8879) );
INV_X32 U_I16150 ( .A(g3900), .ZN(I16150) );
INV_X32 U_g8882 ( .A(I16150), .ZN(g8882) );
INV_X32 U_I16153 ( .A(g3306), .ZN(I16153) );
INV_X32 U_g8885 ( .A(I16153), .ZN(g8885) );
INV_X32 U_I16156 ( .A(g5438), .ZN(I16156) );
INV_X32 U_g8888 ( .A(I16156), .ZN(g8888) );
INV_X32 U_I16159 ( .A(g5403), .ZN(I16159) );
INV_X32 U_g8891 ( .A(I16159), .ZN(g8891) );
INV_X32 U_I16163 ( .A(g6031), .ZN(I16163) );
INV_X32 U_g8893 ( .A(I16163), .ZN(g8893) );
INV_X32 U_I16166 ( .A(g6713), .ZN(I16166) );
INV_X32 U_g8894 ( .A(I16166), .ZN(g8894) );
INV_X32 U_I16169 ( .A(g5405), .ZN(I16169) );
INV_X32 U_g8897 ( .A(I16169), .ZN(g8897) );
INV_X32 U_I16172 ( .A(g5413), .ZN(I16172) );
INV_X32 U_g8898 ( .A(I16172), .ZN(g8898) );
INV_X32 U_I16176 ( .A(g7936), .ZN(I16176) );
INV_X32 U_g8900 ( .A(I16176), .ZN(g8900) );
INV_X32 U_I16179 ( .A(g5512), .ZN(I16179) );
INV_X32 U_g8901 ( .A(I16179), .ZN(g8901) );
INV_X32 U_I16182 ( .A(g5407), .ZN(I16182) );
INV_X32 U_g8904 ( .A(I16182), .ZN(g8904) );
INV_X32 U_I16185 ( .A(g5415), .ZN(I16185) );
INV_X32 U_g8905 ( .A(I16185), .ZN(g8905) );
INV_X32 U_I16190 ( .A(g6118), .ZN(I16190) );
INV_X32 U_g8908 ( .A(I16190), .ZN(g8908) );
INV_X32 U_I16193 ( .A(g5417), .ZN(I16193) );
INV_X32 U_g8909 ( .A(I16193), .ZN(g8909) );
INV_X32 U_I16196 ( .A(g6116), .ZN(I16196) );
INV_X32 U_g8910 ( .A(I16196), .ZN(g8910) );
INV_X32 U_g8911 ( .A(g5114), .ZN(g8911) );
INV_X32 U_I16200 ( .A(g7303), .ZN(I16200) );
INV_X32 U_g8912 ( .A(I16200), .ZN(g8912) );
INV_X32 U_I16203 ( .A(g3878), .ZN(I16203) );
INV_X32 U_g8915 ( .A(I16203), .ZN(g8915) );
INV_X32 U_I16206 ( .A(g6448), .ZN(I16206) );
INV_X32 U_g8918 ( .A(I16206), .ZN(g8918) );
INV_X32 U_I16209 ( .A(g5438), .ZN(I16209) );
INV_X32 U_g8921 ( .A(I16209), .ZN(g8921) );
INV_X32 U_I16212 ( .A(g5411), .ZN(I16212) );
INV_X32 U_g8924 ( .A(I16212), .ZN(g8924) );
INV_X32 U_I16215 ( .A(g3462), .ZN(I16215) );
INV_X32 U_g8925 ( .A(I16215), .ZN(g8925) );
INV_X32 U_I16218 ( .A(g5473), .ZN(I16218) );
INV_X32 U_g8928 ( .A(I16218), .ZN(g8928) );
INV_X32 U_I16221 ( .A(g5412), .ZN(I16221) );
INV_X32 U_g8931 ( .A(I16221), .ZN(g8931) );
INV_X32 U_I16225 ( .A(g6042), .ZN(I16225) );
INV_X32 U_g8933 ( .A(I16225), .ZN(g8933) );
INV_X32 U_I16228 ( .A(g7015), .ZN(I16228) );
INV_X32 U_g8934 ( .A(I16228), .ZN(g8934) );
INV_X32 U_I16231 ( .A(g5414), .ZN(I16231) );
INV_X32 U_g8937 ( .A(I16231), .ZN(g8937) );
INV_X32 U_I16234 ( .A(g5420), .ZN(I16234) );
INV_X32 U_g8938 ( .A(I16234), .ZN(g8938) );
INV_X32 U_I16238 ( .A(g7936), .ZN(I16238) );
INV_X32 U_g8940 ( .A(I16238), .ZN(g8940) );
INV_X32 U_I16241 ( .A(g5556), .ZN(I16241) );
INV_X32 U_g8941 ( .A(I16241), .ZN(g8941) );
INV_X32 U_I16244 ( .A(g5416), .ZN(I16244) );
INV_X32 U_g8944 ( .A(I16244), .ZN(g8944) );
INV_X32 U_I16247 ( .A(g5422), .ZN(I16247) );
INV_X32 U_g8945 ( .A(I16247), .ZN(g8945) );
INV_X32 U_I16252 ( .A(g6134), .ZN(I16252) );
INV_X32 U_g8948 ( .A(I16252), .ZN(g8948) );
INV_X32 U_I16255 ( .A(g3900), .ZN(I16255) );
INV_X32 U_g8949 ( .A(I16255), .ZN(g8949) );
INV_X32 U_I16258 ( .A(g3306), .ZN(I16258) );
INV_X32 U_g8952 ( .A(I16258), .ZN(g8952) );
INV_X32 U_I16261 ( .A(g6448), .ZN(I16261) );
INV_X32 U_g8955 ( .A(I16261), .ZN(g8955) );
INV_X32 U_I16264 ( .A(g6713), .ZN(I16264) );
INV_X32 U_g8958 ( .A(I16264), .ZN(g8958) );
INV_X32 U_I16267 ( .A(g5473), .ZN(I16267) );
INV_X32 U_g8961 ( .A(I16267), .ZN(g8961) );
INV_X32 U_I16270 ( .A(g5418), .ZN(I16270) );
INV_X32 U_g8964 ( .A(I16270), .ZN(g8964) );
INV_X32 U_I16273 ( .A(g3618), .ZN(I16273) );
INV_X32 U_g8965 ( .A(I16273), .ZN(g8965) );
INV_X32 U_I16276 ( .A(g5512), .ZN(I16276) );
INV_X32 U_g8968 ( .A(I16276), .ZN(g8968) );
INV_X32 U_I16279 ( .A(g5419), .ZN(I16279) );
INV_X32 U_g8971 ( .A(I16279), .ZN(g8971) );
INV_X32 U_I16283 ( .A(g6046), .ZN(I16283) );
INV_X32 U_g8973 ( .A(I16283), .ZN(g8973) );
INV_X32 U_I16286 ( .A(g7265), .ZN(I16286) );
INV_X32 U_g8974 ( .A(I16286), .ZN(g8974) );
INV_X32 U_I16289 ( .A(g5421), .ZN(I16289) );
INV_X32 U_g8977 ( .A(I16289), .ZN(g8977) );
INV_X32 U_I16292 ( .A(g5426), .ZN(I16292) );
INV_X32 U_g8978 ( .A(I16292), .ZN(g8978) );
INV_X32 U_I16296 ( .A(g3306), .ZN(I16296) );
INV_X32 U_g8980 ( .A(I16296), .ZN(g8980) );
INV_X32 U_g8983 ( .A(g6486), .ZN(g8983) );
INV_X32 U_I16300 ( .A(g3462), .ZN(I16300) );
INV_X32 U_g8984 ( .A(I16300), .ZN(g8984) );
INV_X32 U_I16303 ( .A(g6713), .ZN(I16303) );
INV_X32 U_g8987 ( .A(I16303), .ZN(g8987) );
INV_X32 U_I16306 ( .A(g7015), .ZN(I16306) );
INV_X32 U_g8990 ( .A(I16306), .ZN(g8990) );
INV_X32 U_I16309 ( .A(g5512), .ZN(I16309) );
INV_X32 U_g8993 ( .A(I16309), .ZN(g8993) );
INV_X32 U_I16312 ( .A(g5424), .ZN(I16312) );
INV_X32 U_g8996 ( .A(I16312), .ZN(g8996) );
INV_X32 U_I16315 ( .A(g3774), .ZN(I16315) );
INV_X32 U_g8997 ( .A(I16315), .ZN(g8997) );
INV_X32 U_I16318 ( .A(g5556), .ZN(I16318) );
INV_X32 U_g9000 ( .A(I16318), .ZN(g9000) );
INV_X32 U_I16321 ( .A(g5425), .ZN(I16321) );
INV_X32 U_g9003 ( .A(I16321), .ZN(g9003) );
INV_X32 U_I16325 ( .A(g6052), .ZN(I16325) );
INV_X32 U_g9005 ( .A(I16325), .ZN(g9005) );
INV_X32 U_I16328 ( .A(g3900), .ZN(I16328) );
INV_X32 U_g9006 ( .A(I16328), .ZN(g9006) );
INV_X32 U_I16332 ( .A(g3462), .ZN(I16332) );
INV_X32 U_g9010 ( .A(I16332), .ZN(g9010) );
INV_X32 U_I16335 ( .A(g3618), .ZN(I16335) );
INV_X32 U_g9013 ( .A(I16335), .ZN(g9013) );
INV_X32 U_I16338 ( .A(g7015), .ZN(I16338) );
INV_X32 U_g9016 ( .A(I16338), .ZN(g9016) );
INV_X32 U_I16341 ( .A(g7265), .ZN(I16341) );
INV_X32 U_g9019 ( .A(I16341), .ZN(g9019) );
INV_X32 U_I16344 ( .A(g5556), .ZN(I16344) );
INV_X32 U_g9022 ( .A(I16344), .ZN(g9022) );
INV_X32 U_I16347 ( .A(g5427), .ZN(I16347) );
INV_X32 U_g9025 ( .A(I16347), .ZN(g9025) );
INV_X32 U_g9027 ( .A(g5679), .ZN(g9027) );
INV_X32 U_I16354 ( .A(g3618), .ZN(I16354) );
INV_X32 U_g9035 ( .A(I16354), .ZN(g9035) );
INV_X32 U_I16357 ( .A(g3774), .ZN(I16357) );
INV_X32 U_g9038 ( .A(I16357), .ZN(g9038) );
INV_X32 U_I16360 ( .A(g7265), .ZN(I16360) );
INV_X32 U_g9041 ( .A(I16360), .ZN(g9041) );
INV_X32 U_I16363 ( .A(g3900), .ZN(I16363) );
INV_X32 U_g9044 ( .A(I16363), .ZN(g9044) );
INV_X32 U_g9050 ( .A(g5731), .ZN(g9050) );
INV_X32 U_I16372 ( .A(g3774), .ZN(I16372) );
INV_X32 U_g9058 ( .A(I16372), .ZN(g9058) );
INV_X32 U_g9067 ( .A(g5789), .ZN(g9067) );
INV_X32 U_g9084 ( .A(g5848), .ZN(g9084) );
INV_X32 U_I16432 ( .A(g3366), .ZN(I16432) );
INV_X32 U_g9128 ( .A(I16432), .ZN(g9128) );
INV_X32 U_I16438 ( .A(g3522), .ZN(I16438) );
INV_X32 U_g9134 ( .A(I16438), .ZN(g9134) );
INV_X32 U_I16444 ( .A(g3678), .ZN(I16444) );
INV_X32 U_g9140 ( .A(I16444), .ZN(g9140) );
INV_X32 U_I16450 ( .A(g3834), .ZN(I16450) );
INV_X32 U_g9146 ( .A(I16450), .ZN(g9146) );
INV_X32 U_I16453 ( .A(g7936), .ZN(I16453) );
INV_X32 U_g9149 ( .A(I16453), .ZN(g9149) );
INV_X32 U_g9150 ( .A(g5893), .ZN(g9150) );
INV_X32 U_I16457 ( .A(g7936), .ZN(I16457) );
INV_X32 U_g9159 ( .A(I16457), .ZN(g9159) );
INV_X32 U_g9160 ( .A(g6170), .ZN(g9160) );
INV_X32 U_g9161 ( .A(g5852), .ZN(g9161) );
INV_X32 U_I16462 ( .A(g5438), .ZN(I16462) );
INV_X32 U_g9170 ( .A(I16462), .ZN(g9170) );
INV_X32 U_I16465 ( .A(g6000), .ZN(I16465) );
INV_X32 U_g9173 ( .A(I16465), .ZN(g9173) );
INV_X32 U_g9174 ( .A(g5932), .ZN(g9174) );
INV_X32 U_I16469 ( .A(g7936), .ZN(I16469) );
INV_X32 U_g9183 ( .A(I16469), .ZN(g9183) );
INV_X32 U_I16472 ( .A(g7901), .ZN(I16472) );
INV_X32 U_g9184 ( .A(I16472), .ZN(g9184) );
INV_X32 U_g9187 ( .A(g5803), .ZN(g9187) );
INV_X32 U_I16476 ( .A(g6448), .ZN(I16476) );
INV_X32 U_g9196 ( .A(I16476), .ZN(g9196) );
INV_X32 U_I16479 ( .A(g5438), .ZN(I16479) );
INV_X32 U_g9199 ( .A(I16479), .ZN(g9199) );
INV_X32 U_I16482 ( .A(g6000), .ZN(I16482) );
INV_X32 U_g9202 ( .A(I16482), .ZN(g9202) );
INV_X32 U_g9203 ( .A(g5899), .ZN(g9203) );
INV_X32 U_I16486 ( .A(g5473), .ZN(I16486) );
INV_X32 U_g9212 ( .A(I16486), .ZN(g9212) );
INV_X32 U_I16489 ( .A(g6000), .ZN(I16489) );
INV_X32 U_g9215 ( .A(I16489), .ZN(g9215) );
INV_X32 U_g9216 ( .A(g5966), .ZN(g9216) );
INV_X32 U_I16493 ( .A(g7936), .ZN(I16493) );
INV_X32 U_g9225 ( .A(I16493), .ZN(g9225) );
INV_X32 U_g9226 ( .A(g5434), .ZN(g9226) );
INV_X32 U_g9227 ( .A(g5587), .ZN(g9227) );
INV_X32 U_g9228 ( .A(g7667), .ZN(g9228) );
INV_X32 U_I16499 ( .A(g7901), .ZN(I16499) );
INV_X32 U_g9229 ( .A(I16499), .ZN(g9229) );
INV_X32 U_g9232 ( .A(g5752), .ZN(g9232) );
INV_X32 U_I16504 ( .A(g3306), .ZN(I16504) );
INV_X32 U_g9242 ( .A(I16504), .ZN(g9242) );
INV_X32 U_I16507 ( .A(g6448), .ZN(I16507) );
INV_X32 U_g9245 ( .A(I16507), .ZN(g9245) );
INV_X32 U_g9248 ( .A(g5859), .ZN(g9248) );
INV_X32 U_I16511 ( .A(g6713), .ZN(I16511) );
INV_X32 U_g9257 ( .A(I16511), .ZN(g9257) );
INV_X32 U_I16514 ( .A(g5473), .ZN(I16514) );
INV_X32 U_g9260 ( .A(I16514), .ZN(g9260) );
INV_X32 U_I16517 ( .A(g6000), .ZN(I16517) );
INV_X32 U_g9263 ( .A(I16517), .ZN(g9263) );
INV_X32 U_g9264 ( .A(g5938), .ZN(g9264) );
INV_X32 U_I16521 ( .A(g5512), .ZN(I16521) );
INV_X32 U_g9273 ( .A(I16521), .ZN(g9273) );
INV_X32 U_I16524 ( .A(g6000), .ZN(I16524) );
INV_X32 U_g9276 ( .A(I16524), .ZN(g9276) );
INV_X32 U_g9277 ( .A(g5995), .ZN(g9277) );
INV_X32 U_g9286 ( .A(g6197), .ZN(g9286) );
INV_X32 U_g9287 ( .A(g6638), .ZN(g9287) );
INV_X32 U_g9288 ( .A(g5363), .ZN(g9288) );
INV_X32 U_g9289 ( .A(g5379), .ZN(g9289) );
INV_X32 U_I16532 ( .A(g7901), .ZN(I16532) );
INV_X32 U_g9290 ( .A(I16532), .ZN(g9290) );
INV_X32 U_g9293 ( .A(g5703), .ZN(g9293) );
INV_X32 U_I16538 ( .A(g3306), .ZN(I16538) );
INV_X32 U_g9303 ( .A(I16538), .ZN(g9303) );
INV_X32 U_I16541 ( .A(g5438), .ZN(I16541) );
INV_X32 U_g9306 ( .A(I16541), .ZN(g9306) );
INV_X32 U_I16544 ( .A(g6054), .ZN(I16544) );
INV_X32 U_g9309 ( .A(I16544), .ZN(g9309) );
INV_X32 U_g9310 ( .A(g5811), .ZN(g9310) );
INV_X32 U_I16549 ( .A(g3462), .ZN(I16549) );
INV_X32 U_g9320 ( .A(I16549), .ZN(g9320) );
INV_X32 U_I16552 ( .A(g6713), .ZN(I16552) );
INV_X32 U_g9323 ( .A(I16552), .ZN(g9323) );
INV_X32 U_g9326 ( .A(g5906), .ZN(g9326) );
INV_X32 U_I16556 ( .A(g7015), .ZN(I16556) );
INV_X32 U_g9335 ( .A(I16556), .ZN(g9335) );
INV_X32 U_I16559 ( .A(g5512), .ZN(I16559) );
INV_X32 U_g9338 ( .A(I16559), .ZN(g9338) );
INV_X32 U_I16562 ( .A(g6000), .ZN(I16562) );
INV_X32 U_g9341 ( .A(I16562), .ZN(g9341) );
INV_X32 U_g9342 ( .A(g5972), .ZN(g9342) );
INV_X32 U_I16566 ( .A(g5556), .ZN(I16566) );
INV_X32 U_g9351 ( .A(I16566), .ZN(g9351) );
INV_X32 U_I16569 ( .A(g6000), .ZN(I16569) );
INV_X32 U_g9354 ( .A(I16569), .ZN(g9354) );
INV_X32 U_g9355 ( .A(g7639), .ZN(g9355) );
INV_X32 U_g9356 ( .A(g5665), .ZN(g9356) );
INV_X32 U_I16578 ( .A(g6448), .ZN(I16578) );
INV_X32 U_g9368 ( .A(I16578), .ZN(g9368) );
INV_X32 U_I16581 ( .A(g5438), .ZN(I16581) );
INV_X32 U_g9371 ( .A(I16581), .ZN(g9371) );
INV_X32 U_g9374 ( .A(g5761), .ZN(g9374) );
INV_X32 U_I16587 ( .A(g3462), .ZN(I16587) );
INV_X32 U_g9384 ( .A(I16587), .ZN(g9384) );
INV_X32 U_I16590 ( .A(g5473), .ZN(I16590) );
INV_X32 U_g9387 ( .A(I16590), .ZN(g9387) );
INV_X32 U_I16593 ( .A(g6059), .ZN(I16593) );
INV_X32 U_g9390 ( .A(I16593), .ZN(g9390) );
INV_X32 U_g9391 ( .A(g5867), .ZN(g9391) );
INV_X32 U_I16598 ( .A(g3618), .ZN(I16598) );
INV_X32 U_g9401 ( .A(I16598), .ZN(g9401) );
INV_X32 U_I16601 ( .A(g7015), .ZN(I16601) );
INV_X32 U_g9404 ( .A(I16601), .ZN(g9404) );
INV_X32 U_g9407 ( .A(g5945), .ZN(g9407) );
INV_X32 U_I16605 ( .A(g7265), .ZN(I16605) );
INV_X32 U_g9416 ( .A(I16605), .ZN(g9416) );
INV_X32 U_I16608 ( .A(g5556), .ZN(I16608) );
INV_X32 U_g9419 ( .A(I16608), .ZN(g9419) );
INV_X32 U_I16611 ( .A(g6000), .ZN(I16611) );
INV_X32 U_g9422 ( .A(I16611), .ZN(g9422) );
INV_X32 U_g9423 ( .A(g5428), .ZN(g9423) );
INV_X32 U_g9424 ( .A(g5469), .ZN(g9424) );
INV_X32 U_g9425 ( .A(g5346), .ZN(g9425) );
INV_X32 U_g9426 ( .A(g5543), .ZN(g9426) );
INV_X32 U_g9427 ( .A(g5645), .ZN(g9427) );
INV_X32 U_I16624 ( .A(g3306), .ZN(I16624) );
INV_X32 U_g9443 ( .A(I16624), .ZN(g9443) );
INV_X32 U_I16627 ( .A(g6448), .ZN(I16627) );
INV_X32 U_g9446 ( .A(I16627), .ZN(g9446) );
INV_X32 U_I16630 ( .A(g6057), .ZN(I16630) );
INV_X32 U_g9449 ( .A(I16630), .ZN(g9449) );
INV_X32 U_I16633 ( .A(g6486), .ZN(I16633) );
INV_X32 U_g9450 ( .A(I16633), .ZN(g9450) );
INV_X32 U_g9453 ( .A(g5717), .ZN(g9453) );
INV_X32 U_I16641 ( .A(g6713), .ZN(I16641) );
INV_X32 U_g9465 ( .A(I16641), .ZN(g9465) );
INV_X32 U_I16644 ( .A(g5473), .ZN(I16644) );
INV_X32 U_g9468 ( .A(I16644), .ZN(g9468) );
INV_X32 U_g9471 ( .A(g5820), .ZN(g9471) );
INV_X32 U_I16650 ( .A(g3618), .ZN(I16650) );
INV_X32 U_g9481 ( .A(I16650), .ZN(g9481) );
INV_X32 U_I16653 ( .A(g5512), .ZN(I16653) );
INV_X32 U_g9484 ( .A(I16653), .ZN(g9484) );
INV_X32 U_I16656 ( .A(g6066), .ZN(I16656) );
INV_X32 U_g9487 ( .A(I16656), .ZN(g9487) );
INV_X32 U_g9488 ( .A(g5914), .ZN(g9488) );
INV_X32 U_I16661 ( .A(g3774), .ZN(I16661) );
INV_X32 U_g9498 ( .A(I16661), .ZN(g9498) );
INV_X32 U_I16664 ( .A(g7265), .ZN(I16664) );
INV_X32 U_g9501 ( .A(I16664), .ZN(g9501) );
INV_X32 U_g9504 ( .A(g6149), .ZN(g9504) );
INV_X32 U_g9505 ( .A(g6227), .ZN(g9505) );
INV_X32 U_g9506 ( .A(g6444), .ZN(g9506) );
INV_X32 U_g9507 ( .A(g5953), .ZN(g9507) );
INV_X32 U_I16677 ( .A(g3306), .ZN(I16677) );
INV_X32 U_g9524 ( .A(I16677), .ZN(g9524) );
INV_X32 U_g9527 ( .A(g5508), .ZN(g9527) );
INV_X32 U_I16681 ( .A(g6643), .ZN(I16681) );
INV_X32 U_g9528 ( .A(I16681), .ZN(g9528) );
INV_X32 U_I16684 ( .A(g6486), .ZN(I16684) );
INV_X32 U_g9531 ( .A(I16684), .ZN(g9531) );
INV_X32 U_g9569 ( .A(g5683), .ZN(g9569) );
INV_X32 U_I16694 ( .A(g3462), .ZN(I16694) );
INV_X32 U_g9585 ( .A(I16694), .ZN(g9585) );
INV_X32 U_I16697 ( .A(g6713), .ZN(I16697) );
INV_X32 U_g9588 ( .A(I16697), .ZN(g9588) );
INV_X32 U_I16700 ( .A(g6064), .ZN(I16700) );
INV_X32 U_g9591 ( .A(I16700), .ZN(g9591) );
INV_X32 U_I16703 ( .A(g6751), .ZN(I16703) );
INV_X32 U_g9592 ( .A(I16703), .ZN(g9592) );
INV_X32 U_g9595 ( .A(g5775), .ZN(g9595) );
INV_X32 U_I16711 ( .A(g7015), .ZN(I16711) );
INV_X32 U_g9607 ( .A(I16711), .ZN(g9607) );
INV_X32 U_I16714 ( .A(g5512), .ZN(I16714) );
INV_X32 U_g9610 ( .A(I16714), .ZN(g9610) );
INV_X32 U_g9613 ( .A(g5876), .ZN(g9613) );
INV_X32 U_I16720 ( .A(g3774), .ZN(I16720) );
INV_X32 U_g9623 ( .A(I16720), .ZN(g9623) );
INV_X32 U_I16723 ( .A(g5556), .ZN(I16723) );
INV_X32 U_g9626 ( .A(I16723), .ZN(g9626) );
INV_X32 U_I16726 ( .A(g6085), .ZN(I16726) );
INV_X32 U_g9629 ( .A(I16726), .ZN(g9629) );
INV_X32 U_I16741 ( .A(g6062), .ZN(I16741) );
INV_X32 U_g9640 ( .A(I16741), .ZN(g9640) );
INV_X32 U_I16744 ( .A(g3338), .ZN(I16744) );
INV_X32 U_g9641 ( .A(I16744), .ZN(g9641) );
INV_X32 U_I16747 ( .A(g6643), .ZN(I16747) );
INV_X32 U_g9644 ( .A(I16747), .ZN(g9644) );
INV_X32 U_g9649 ( .A(g5982), .ZN(g9649) );
INV_X32 U_I16759 ( .A(g3462), .ZN(I16759) );
INV_X32 U_g9666 ( .A(I16759), .ZN(g9666) );
INV_X32 U_g9669 ( .A(g5552), .ZN(g9669) );
INV_X32 U_I16763 ( .A(g6945), .ZN(I16763) );
INV_X32 U_g9670 ( .A(I16763), .ZN(g9670) );
INV_X32 U_I16766 ( .A(g6751), .ZN(I16766) );
INV_X32 U_g9673 ( .A(I16766), .ZN(g9673) );
INV_X32 U_g9711 ( .A(g5735), .ZN(g9711) );
INV_X32 U_I16776 ( .A(g3618), .ZN(I16776) );
INV_X32 U_g9727 ( .A(I16776), .ZN(g9727) );
INV_X32 U_I16779 ( .A(g7015), .ZN(I16779) );
INV_X32 U_g9730 ( .A(I16779), .ZN(g9730) );
INV_X32 U_I16782 ( .A(g6083), .ZN(I16782) );
INV_X32 U_g9733 ( .A(I16782), .ZN(g9733) );
INV_X32 U_I16785 ( .A(g7053), .ZN(I16785) );
INV_X32 U_g9734 ( .A(I16785), .ZN(g9734) );
INV_X32 U_g9737 ( .A(g5834), .ZN(g9737) );
INV_X32 U_I16793 ( .A(g7265), .ZN(I16793) );
INV_X32 U_g9749 ( .A(I16793), .ZN(g9749) );
INV_X32 U_I16796 ( .A(g5556), .ZN(I16796) );
INV_X32 U_g9752 ( .A(I16796), .ZN(g9752) );
INV_X32 U_g9755 ( .A(g5431), .ZN(g9755) );
INV_X32 U_g9756 ( .A(g5504), .ZN(g9756) );
INV_X32 U_g9757 ( .A(g5601), .ZN(g9757) );
INV_X32 U_g9758 ( .A(g5618), .ZN(g9758) );
INV_X32 U_I16811 ( .A(g3338), .ZN(I16811) );
INV_X32 U_g9767 ( .A(I16811), .ZN(g9767) );
INV_X32 U_I16814 ( .A(g6486), .ZN(I16814) );
INV_X32 U_g9770 ( .A(I16814), .ZN(g9770) );
INV_X32 U_I16832 ( .A(g6081), .ZN(I16832) );
INV_X32 U_g9786 ( .A(I16832), .ZN(g9786) );
INV_X32 U_I16835 ( .A(g3494), .ZN(I16835) );
INV_X32 U_g9787 ( .A(I16835), .ZN(g9787) );
INV_X32 U_I16838 ( .A(g6945), .ZN(I16838) );
INV_X32 U_g9790 ( .A(I16838), .ZN(g9790) );
INV_X32 U_g9795 ( .A(g6019), .ZN(g9795) );
INV_X32 U_I16850 ( .A(g3618), .ZN(I16850) );
INV_X32 U_g9812 ( .A(I16850), .ZN(g9812) );
INV_X32 U_g9815 ( .A(g5598), .ZN(g9815) );
INV_X32 U_I16854 ( .A(g7195), .ZN(I16854) );
INV_X32 U_g9816 ( .A(I16854), .ZN(g9816) );
INV_X32 U_I16857 ( .A(g7053), .ZN(I16857) );
INV_X32 U_g9819 ( .A(I16857), .ZN(g9819) );
INV_X32 U_g9857 ( .A(g5793), .ZN(g9857) );
INV_X32 U_I16867 ( .A(g3774), .ZN(I16867) );
INV_X32 U_g9873 ( .A(I16867), .ZN(g9873) );
INV_X32 U_I16870 ( .A(g7265), .ZN(I16870) );
INV_X32 U_g9876 ( .A(I16870), .ZN(g9876) );
INV_X32 U_I16873 ( .A(g6102), .ZN(I16873) );
INV_X32 U_g9879 ( .A(I16873), .ZN(g9879) );
INV_X32 U_I16876 ( .A(g7303), .ZN(I16876) );
INV_X32 U_g9880 ( .A(I16876), .ZN(g9880) );
INV_X32 U_g9884 ( .A(g6310), .ZN(g9884) );
INV_X32 U_g9885 ( .A(g6905), .ZN(g9885) );
INV_X32 U_g9886 ( .A(g7149), .ZN(g9886) );
INV_X32 U_I16897 ( .A(g6643), .ZN(I16897) );
INV_X32 U_g9895 ( .A(I16897), .ZN(g9895) );
INV_X32 U_I16900 ( .A(g6486), .ZN(I16900) );
INV_X32 U_g9898 ( .A(I16900), .ZN(g9898) );
INV_X32 U_I16915 ( .A(g3494), .ZN(I16915) );
INV_X32 U_g9913 ( .A(I16915), .ZN(g9913) );
INV_X32 U_I16918 ( .A(g6751), .ZN(I16918) );
INV_X32 U_g9916 ( .A(I16918), .ZN(g9916) );
INV_X32 U_I16936 ( .A(g6100), .ZN(I16936) );
INV_X32 U_g9932 ( .A(I16936), .ZN(g9932) );
INV_X32 U_I16939 ( .A(g3650), .ZN(I16939) );
INV_X32 U_g9933 ( .A(I16939), .ZN(g9933) );
INV_X32 U_I16942 ( .A(g7195), .ZN(I16942) );
INV_X32 U_g9936 ( .A(I16942), .ZN(g9936) );
INV_X32 U_g9941 ( .A(g6035), .ZN(g9941) );
INV_X32 U_I16954 ( .A(g3774), .ZN(I16954) );
INV_X32 U_g9958 ( .A(I16954), .ZN(g9958) );
INV_X32 U_g9961 ( .A(g5615), .ZN(g9961) );
INV_X32 U_I16958 ( .A(g7391), .ZN(I16958) );
INV_X32 U_g9962 ( .A(I16958), .ZN(g9962) );
INV_X32 U_I16961 ( .A(g7303), .ZN(I16961) );
INV_X32 U_g9965 ( .A(I16961), .ZN(g9965) );
INV_X32 U_I16972 ( .A(g3900), .ZN(I16972) );
INV_X32 U_g10004 ( .A(I16972), .ZN(g10004) );
INV_X32 U_g10015 ( .A(g5292), .ZN(g10015) );
INV_X32 U_I16984 ( .A(g7936), .ZN(I16984) );
INV_X32 U_g10016 ( .A(I16984), .ZN(g10016) );
INV_X32 U_I16987 ( .A(g6079), .ZN(I16987) );
INV_X32 U_g10017 ( .A(I16987), .ZN(g10017) );
INV_X32 U_I16990 ( .A(g3338), .ZN(I16990) );
INV_X32 U_g10018 ( .A(I16990), .ZN(g10018) );
INV_X32 U_I16993 ( .A(g6643), .ZN(I16993) );
INV_X32 U_g10021 ( .A(I16993), .ZN(g10021) );
INV_X32 U_I17009 ( .A(g6945), .ZN(I17009) );
INV_X32 U_g10049 ( .A(I17009), .ZN(g10049) );
INV_X32 U_I17012 ( .A(g6751), .ZN(I17012) );
INV_X32 U_g10052 ( .A(I17012), .ZN(g10052) );
INV_X32 U_I17027 ( .A(g3650), .ZN(I17027) );
INV_X32 U_g10067 ( .A(I17027), .ZN(g10067) );
INV_X32 U_I17030 ( .A(g7053), .ZN(I17030) );
INV_X32 U_g10070 ( .A(I17030), .ZN(g10070) );
INV_X32 U_I17048 ( .A(g6117), .ZN(I17048) );
INV_X32 U_g10086 ( .A(I17048), .ZN(g10086) );
INV_X32 U_I17051 ( .A(g3806), .ZN(I17051) );
INV_X32 U_g10087 ( .A(I17051), .ZN(g10087) );
INV_X32 U_I17054 ( .A(g7391), .ZN(I17054) );
INV_X32 U_g10090 ( .A(I17054), .ZN(g10090) );
INV_X32 U_I17066 ( .A(g3900), .ZN(I17066) );
INV_X32 U_g10096 ( .A(I17066), .ZN(g10096) );
INV_X32 U_g10099 ( .A(g7700), .ZN(g10099) );
INV_X32 U_I17070 ( .A(g7528), .ZN(I17070) );
INV_X32 U_g10100 ( .A(I17070), .ZN(g10100) );
INV_X32 U_I17081 ( .A(g3338), .ZN(I17081) );
INV_X32 U_g10109 ( .A(I17081), .ZN(g10109) );
INV_X32 U_g10124 ( .A(g5326), .ZN(g10124) );
INV_X32 U_I17097 ( .A(g7936), .ZN(I17097) );
INV_X32 U_g10125 ( .A(I17097), .ZN(g10125) );
INV_X32 U_I17100 ( .A(g6098), .ZN(I17100) );
INV_X32 U_g10126 ( .A(I17100), .ZN(g10126) );
INV_X32 U_I17103 ( .A(g3494), .ZN(I17103) );
INV_X32 U_g10127 ( .A(I17103), .ZN(g10127) );
INV_X32 U_I17106 ( .A(g6945), .ZN(I17106) );
INV_X32 U_g10130 ( .A(I17106), .ZN(g10130) );
INV_X32 U_I17122 ( .A(g7195), .ZN(I17122) );
INV_X32 U_g10158 ( .A(I17122), .ZN(g10158) );
INV_X32 U_I17125 ( .A(g7053), .ZN(I17125) );
INV_X32 U_g10161 ( .A(I17125), .ZN(g10161) );
INV_X32 U_I17140 ( .A(g3806), .ZN(I17140) );
INV_X32 U_g10176 ( .A(I17140), .ZN(g10176) );
INV_X32 U_I17143 ( .A(g7303), .ZN(I17143) );
INV_X32 U_g10179 ( .A(I17143), .ZN(g10179) );
INV_X32 U_I17159 ( .A(g3900), .ZN(I17159) );
INV_X32 U_g10189 ( .A(I17159), .ZN(g10189) );
INV_X32 U_I17184 ( .A(g3494), .ZN(I17184) );
INV_X32 U_g10214 ( .A(I17184), .ZN(g10214) );
INV_X32 U_g10229 ( .A(g5349), .ZN(g10229) );
INV_X32 U_I17200 ( .A(g7936), .ZN(I17200) );
INV_X32 U_g10230 ( .A(I17200), .ZN(g10230) );
INV_X32 U_I17203 ( .A(g6115), .ZN(I17203) );
INV_X32 U_g10231 ( .A(I17203), .ZN(g10231) );
INV_X32 U_I17206 ( .A(g3650), .ZN(I17206) );
INV_X32 U_g10232 ( .A(I17206), .ZN(g10232) );
INV_X32 U_I17209 ( .A(g7195), .ZN(I17209) );
INV_X32 U_g10235 ( .A(I17209), .ZN(g10235) );
INV_X32 U_I17225 ( .A(g7391), .ZN(I17225) );
INV_X32 U_g10263 ( .A(I17225), .ZN(g10263) );
INV_X32 U_I17228 ( .A(g7303), .ZN(I17228) );
INV_X32 U_g10266 ( .A(I17228), .ZN(g10266) );
INV_X32 U_I17235 ( .A(g3900), .ZN(I17235) );
INV_X32 U_g10273 ( .A(I17235), .ZN(g10273) );
INV_X32 U_I17238 ( .A(g3900), .ZN(I17238) );
INV_X32 U_g10276 ( .A(I17238), .ZN(g10276) );
INV_X32 U_I17278 ( .A(g3650), .ZN(I17278) );
INV_X32 U_g10316 ( .A(I17278), .ZN(g10316) );
INV_X32 U_g10331 ( .A(g5366), .ZN(g10331) );
INV_X32 U_I17294 ( .A(g7936), .ZN(I17294) );
INV_X32 U_g10332 ( .A(I17294), .ZN(g10332) );
INV_X32 U_I17297 ( .A(g6130), .ZN(I17297) );
INV_X32 U_g10333 ( .A(I17297), .ZN(g10333) );
INV_X32 U_I17300 ( .A(g3806), .ZN(I17300) );
INV_X32 U_g10334 ( .A(I17300), .ZN(g10334) );
INV_X32 U_I17303 ( .A(g7391), .ZN(I17303) );
INV_X32 U_g10337 ( .A(I17303), .ZN(g10337) );
INV_X32 U_I17311 ( .A(g3900), .ZN(I17311) );
INV_X32 U_g10357 ( .A(I17311), .ZN(g10357) );
INV_X32 U_I17363 ( .A(g3806), .ZN(I17363) );
INV_X32 U_g10409 ( .A(I17363), .ZN(g10409) );
INV_X32 U_I17370 ( .A(g3900), .ZN(I17370) );
INV_X32 U_g10416 ( .A(I17370), .ZN(g10416) );
INV_X32 U_I17373 ( .A(g3900), .ZN(I17373) );
INV_X32 U_g10419 ( .A(I17373), .ZN(g10419) );
INV_X32 U_g10424 ( .A(g7910), .ZN(g10424) );
INV_X32 U_g10481 ( .A(g7826), .ZN(g10481) );
INV_X32 U_I17433 ( .A(g3900), .ZN(I17433) );
INV_X32 U_g10482 ( .A(I17433), .ZN(g10482) );
INV_X32 U_g10486 ( .A(g7957), .ZN(g10486) );
INV_X32 U_g10500 ( .A(g7962), .ZN(g10500) );
INV_X32 U_I17483 ( .A(g3900), .ZN(I17483) );
INV_X32 U_g10542 ( .A(I17483), .ZN(g10542) );
INV_X32 U_I17486 ( .A(g3900), .ZN(I17486) );
INV_X32 U_g10545 ( .A(I17486), .ZN(g10545) );
INV_X32 U_g10549 ( .A(g7999), .ZN(g10549) );
INV_X32 U_g10560 ( .A(g8008), .ZN(g10560) );
INV_X32 U_g10574 ( .A(g8013), .ZN(g10574) );
INV_X32 U_I17527 ( .A(g3900), .ZN(I17527) );
INV_X32 U_g10601 ( .A(I17527), .ZN(g10601) );
INV_X32 U_g10606 ( .A(g8074), .ZN(g10606) );
INV_X32 U_g10617 ( .A(g8083), .ZN(g10617) );
INV_X32 U_g10631 ( .A(g8088), .ZN(g10631) );
INV_X32 U_I17557 ( .A(g3900), .ZN(I17557) );
INV_X32 U_g10646 ( .A(I17557), .ZN(g10646) );
INV_X32 U_g10653 ( .A(g8159), .ZN(g10653) );
INV_X32 U_g10664 ( .A(g8168), .ZN(g10664) );
INV_X32 U_g10683 ( .A(g8245), .ZN(g10683) );
INV_X32 U_g10694 ( .A(g4326), .ZN(g10694) );
INV_X32 U_g10714 ( .A(g4495), .ZN(g10714) );
INV_X32 U_g10730 ( .A(g6173), .ZN(g10730) );
INV_X32 U_g10735 ( .A(g4671), .ZN(g10735) );
INV_X32 U_g10749 ( .A(g6205), .ZN(g10749) );
INV_X32 U_g10754 ( .A(g4848), .ZN(g10754) );
INV_X32 U_g10765 ( .A(g6048), .ZN(g10765) );
INV_X32 U_g10766 ( .A(g6676), .ZN(g10766) );
INV_X32 U_g10767 ( .A(g6294), .ZN(g10767) );
INV_X32 U_g10772 ( .A(g6978), .ZN(g10772) );
INV_X32 U_g10773 ( .A(g6431), .ZN(g10773) );
INV_X32 U_I17627 ( .A(g7575), .ZN(I17627) );
INV_X32 U_g10779 ( .A(I17627), .ZN(g10779) );
INV_X32 U_g10783 ( .A(g7228), .ZN(g10783) );
INV_X32 U_I17632 ( .A(g6183), .ZN(I17632) );
INV_X32 U_g10787 ( .A(I17632), .ZN(g10787) );
INV_X32 U_g10788 ( .A(g7424), .ZN(g10788) );
INV_X32 U_I17637 ( .A(g6204), .ZN(I17637) );
INV_X32 U_g10792 ( .A(I17637), .ZN(g10792) );
INV_X32 U_I17641 ( .A(g6215), .ZN(I17641) );
INV_X32 U_g10796 ( .A(I17641), .ZN(g10796) );
INV_X32 U_I17645 ( .A(g6288), .ZN(I17645) );
INV_X32 U_g10800 ( .A(I17645), .ZN(g10800) );
INV_X32 U_I17649 ( .A(g6293), .ZN(I17649) );
INV_X32 U_g10804 ( .A(I17649), .ZN(g10804) );
INV_X32 U_I17653 ( .A(g6304), .ZN(I17653) );
INV_X32 U_g10808 ( .A(I17653), .ZN(g10808) );
INV_X32 U_g10809 ( .A(g5701), .ZN(g10809) );
INV_X32 U_I17658 ( .A(g6367), .ZN(I17658) );
INV_X32 U_g10813 ( .A(I17658), .ZN(g10813) );
INV_X32 U_I17662 ( .A(g6425), .ZN(I17662) );
INV_X32 U_g10817 ( .A(I17662), .ZN(g10817) );
INV_X32 U_I17666 ( .A(g6430), .ZN(I17666) );
INV_X32 U_g10821 ( .A(I17666), .ZN(g10821) );
INV_X32 U_I17670 ( .A(g6441), .ZN(I17670) );
INV_X32 U_g10825 ( .A(I17670), .ZN(g10825) );
INV_X32 U_I17673 ( .A(g8107), .ZN(I17673) );
INV_X32 U_g10826 ( .A(I17673), .ZN(g10826) );
INV_X32 U_g10829 ( .A(g5749), .ZN(g10829) );
INV_X32 U_I17677 ( .A(g6517), .ZN(I17677) );
INV_X32 U_g10830 ( .A(I17677), .ZN(g10830) );
INV_X32 U_I17681 ( .A(g6572), .ZN(I17681) );
INV_X32 U_g10834 ( .A(I17681), .ZN(g10834) );
INV_X32 U_I17685 ( .A(g6630), .ZN(I17685) );
INV_X32 U_g10838 ( .A(I17685), .ZN(g10838) );
INV_X32 U_I17689 ( .A(g6635), .ZN(I17689) );
INV_X32 U_g10842 ( .A(I17689), .ZN(g10842) );
INV_X32 U_I17692 ( .A(g8107), .ZN(I17692) );
INV_X32 U_g10843 ( .A(I17692), .ZN(g10843) );
INV_X32 U_g10846 ( .A(g5799), .ZN(g10846) );
INV_X32 U_g10847 ( .A(g5800), .ZN(g10847) );
INV_X32 U_g10848 ( .A(g5801), .ZN(g10848) );
INV_X32 U_I17698 ( .A(g6711), .ZN(I17698) );
INV_X32 U_g10849 ( .A(I17698), .ZN(g10849) );
INV_X32 U_I17701 ( .A(g6781), .ZN(I17701) );
INV_X32 U_g10850 ( .A(I17701), .ZN(g10850) );
INV_X32 U_I17705 ( .A(g6836), .ZN(I17705) );
INV_X32 U_g10854 ( .A(I17705), .ZN(g10854) );
INV_X32 U_I17709 ( .A(g6894), .ZN(I17709) );
INV_X32 U_g10858 ( .A(I17709), .ZN(g10858) );
INV_X32 U_I17712 ( .A(g8031), .ZN(I17712) );
INV_X32 U_g10859 ( .A(I17712), .ZN(g10859) );
INV_X32 U_I17715 ( .A(g8107), .ZN(I17715) );
INV_X32 U_g10862 ( .A(I17715), .ZN(g10862) );
INV_X32 U_g10865 ( .A(g6131), .ZN(g10865) );
INV_X32 U_g10866 ( .A(g5849), .ZN(g10866) );
INV_X32 U_g10867 ( .A(g5850), .ZN(g10867) );
INV_X32 U_I17721 ( .A(g6641), .ZN(I17721) );
INV_X32 U_g10868 ( .A(I17721), .ZN(g10868) );
INV_X32 U_I17724 ( .A(g6942), .ZN(I17724) );
INV_X32 U_g10869 ( .A(I17724), .ZN(g10869) );
INV_X32 U_I17727 ( .A(g7013), .ZN(I17727) );
INV_X32 U_g10870 ( .A(I17727), .ZN(g10870) );
INV_X32 U_I17730 ( .A(g7083), .ZN(I17730) );
INV_X32 U_g10871 ( .A(I17730), .ZN(g10871) );
INV_X32 U_I17734 ( .A(g7138), .ZN(I17734) );
INV_X32 U_g10875 ( .A(I17734), .ZN(g10875) );
INV_X32 U_I17737 ( .A(g6000), .ZN(I17737) );
INV_X32 U_g10876 ( .A(I17737), .ZN(g10876) );
INV_X32 U_I17740 ( .A(g8031), .ZN(I17740) );
INV_X32 U_g10877 ( .A(I17740), .ZN(g10877) );
INV_X32 U_I17743 ( .A(g8107), .ZN(I17743) );
INV_X32 U_g10880 ( .A(I17743), .ZN(g10880) );
INV_X32 U_I17746 ( .A(g8107), .ZN(I17746) );
INV_X32 U_g10883 ( .A(I17746), .ZN(g10883) );
INV_X32 U_g10886 ( .A(g5889), .ZN(g10886) );
INV_X32 U_I17750 ( .A(g7157), .ZN(I17750) );
INV_X32 U_g10887 ( .A(I17750), .ZN(g10887) );
INV_X32 U_I17753 ( .A(g6943), .ZN(I17753) );
INV_X32 U_g10888 ( .A(I17753), .ZN(g10888) );
INV_X32 U_I17756 ( .A(g7192), .ZN(I17756) );
INV_X32 U_g10889 ( .A(I17756), .ZN(g10889) );
INV_X32 U_I17759 ( .A(g7263), .ZN(I17759) );
INV_X32 U_g10890 ( .A(I17759), .ZN(g10890) );
INV_X32 U_I17762 ( .A(g7333), .ZN(I17762) );
INV_X32 U_g10891 ( .A(I17762), .ZN(g10891) );
INV_X32 U_I17765 ( .A(g7976), .ZN(I17765) );
INV_X32 U_g10892 ( .A(I17765), .ZN(g10892) );
INV_X32 U_I17768 ( .A(g8031), .ZN(I17768) );
INV_X32 U_g10895 ( .A(I17768), .ZN(g10895) );
INV_X32 U_I17771 ( .A(g8107), .ZN(I17771) );
INV_X32 U_g10898 ( .A(I17771), .ZN(g10898) );
INV_X32 U_I17774 ( .A(g8107), .ZN(I17774) );
INV_X32 U_g10901 ( .A(I17774), .ZN(g10901) );
INV_X32 U_g10904 ( .A(g5922), .ZN(g10904) );
INV_X32 U_g10905 ( .A(g5923), .ZN(g10905) );
INV_X32 U_g10906 ( .A(g5924), .ZN(g10906) );
INV_X32 U_I17780 ( .A(g7348), .ZN(I17780) );
INV_X32 U_g10907 ( .A(I17780), .ZN(g10907) );
INV_X32 U_I17783 ( .A(g7353), .ZN(I17783) );
INV_X32 U_g10908 ( .A(I17783), .ZN(g10908) );
INV_X32 U_I17786 ( .A(g7193), .ZN(I17786) );
INV_X32 U_g10909 ( .A(I17786), .ZN(g10909) );
INV_X32 U_I17789 ( .A(g7388), .ZN(I17789) );
INV_X32 U_g10910 ( .A(I17789), .ZN(g10910) );
INV_X32 U_I17792 ( .A(g7459), .ZN(I17792) );
INV_X32 U_g10911 ( .A(I17792), .ZN(g10911) );
INV_X32 U_I17795 ( .A(g7976), .ZN(I17795) );
INV_X32 U_g10912 ( .A(I17795), .ZN(g10912) );
INV_X32 U_I17798 ( .A(g8031), .ZN(I17798) );
INV_X32 U_g10915 ( .A(I17798), .ZN(g10915) );
INV_X32 U_I17801 ( .A(g8107), .ZN(I17801) );
INV_X32 U_g10918 ( .A(I17801), .ZN(g10918) );
INV_X32 U_I17804 ( .A(g8031), .ZN(I17804) );
INV_X32 U_g10921 ( .A(I17804), .ZN(g10921) );
INV_X32 U_I17807 ( .A(g8107), .ZN(I17807) );
INV_X32 U_g10924 ( .A(I17807), .ZN(g10924) );
INV_X32 U_g10927 ( .A(g6153), .ZN(g10927) );
INV_X32 U_g10928 ( .A(g5951), .ZN(g10928) );
INV_X32 U_g10929 ( .A(g5952), .ZN(g10929) );
INV_X32 U_I17813 ( .A(g5707), .ZN(I17813) );
INV_X32 U_g10930 ( .A(I17813), .ZN(g10930) );
INV_X32 U_I17816 ( .A(g7346), .ZN(I17816) );
INV_X32 U_g10931 ( .A(I17816), .ZN(g10931) );
INV_X32 U_I17819 ( .A(g6448), .ZN(I17819) );
INV_X32 U_g10932 ( .A(I17819), .ZN(g10932) );
INV_X32 U_I17822 ( .A(g7478), .ZN(I17822) );
INV_X32 U_g10933 ( .A(I17822), .ZN(g10933) );
INV_X32 U_I17825 ( .A(g7483), .ZN(I17825) );
INV_X32 U_g10934 ( .A(I17825), .ZN(g10934) );
INV_X32 U_I17828 ( .A(g7389), .ZN(I17828) );
INV_X32 U_g10935 ( .A(I17828), .ZN(g10935) );
INV_X32 U_I17831 ( .A(g7518), .ZN(I17831) );
INV_X32 U_g10936 ( .A(I17831), .ZN(g10936) );
INV_X32 U_I17834 ( .A(g7976), .ZN(I17834) );
INV_X32 U_g10937 ( .A(I17834), .ZN(g10937) );
INV_X32 U_I17837 ( .A(g8031), .ZN(I17837) );
INV_X32 U_g10940 ( .A(I17837), .ZN(g10940) );
INV_X32 U_I17840 ( .A(g8107), .ZN(I17840) );
INV_X32 U_g10943 ( .A(I17840), .ZN(g10943) );
INV_X32 U_I17843 ( .A(g8031), .ZN(I17843) );
INV_X32 U_g10946 ( .A(I17843), .ZN(g10946) );
INV_X32 U_I17846 ( .A(g8107), .ZN(I17846) );
INV_X32 U_g10949 ( .A(I17846), .ZN(g10949) );
INV_X32 U_I17849 ( .A(g8103), .ZN(I17849) );
INV_X32 U_g10952 ( .A(I17849), .ZN(g10952) );
INV_X32 U_g10961 ( .A(g5978), .ZN(g10961) );
INV_X32 U_g10962 ( .A(g5979), .ZN(g10962) );
INV_X32 U_I17854 ( .A(g6232), .ZN(I17854) );
INV_X32 U_g10963 ( .A(I17854), .ZN(g10963) );
INV_X32 U_I17857 ( .A(g6448), .ZN(I17857) );
INV_X32 U_g10966 ( .A(I17857), .ZN(g10966) );
INV_X32 U_I17860 ( .A(g5765), .ZN(I17860) );
INV_X32 U_g10967 ( .A(I17860), .ZN(g10967) );
INV_X32 U_I17863 ( .A(g7476), .ZN(I17863) );
INV_X32 U_g10968 ( .A(I17863), .ZN(g10968) );
INV_X32 U_I17866 ( .A(g6713), .ZN(I17866) );
INV_X32 U_g10969 ( .A(I17866), .ZN(g10969) );
INV_X32 U_I17869 ( .A(g7534), .ZN(I17869) );
INV_X32 U_g10972 ( .A(I17869), .ZN(g10972) );
INV_X32 U_I17872 ( .A(g7539), .ZN(I17872) );
INV_X32 U_g10973 ( .A(I17872), .ZN(g10973) );
INV_X32 U_I17875 ( .A(g7976), .ZN(I17875) );
INV_X32 U_g10974 ( .A(I17875), .ZN(g10974) );
INV_X32 U_I17878 ( .A(g8031), .ZN(I17878) );
INV_X32 U_g10977 ( .A(I17878), .ZN(g10977) );
INV_X32 U_I17881 ( .A(g7976), .ZN(I17881) );
INV_X32 U_g10980 ( .A(I17881), .ZN(g10980) );
INV_X32 U_I17884 ( .A(g8031), .ZN(I17884) );
INV_X32 U_g10983 ( .A(I17884), .ZN(g10983) );
INV_X32 U_g10986 ( .A(g6014), .ZN(g10986) );
INV_X32 U_g10987 ( .A(g6015), .ZN(g10987) );
INV_X32 U_I17889 ( .A(g6314), .ZN(I17889) );
INV_X32 U_g10988 ( .A(I17889), .ZN(g10988) );
INV_X32 U_I17892 ( .A(g6232), .ZN(I17892) );
INV_X32 U_g10991 ( .A(I17892), .ZN(g10991) );
INV_X32 U_I17895 ( .A(g6448), .ZN(I17895) );
INV_X32 U_g10994 ( .A(I17895), .ZN(g10994) );
INV_X32 U_I17898 ( .A(g6643), .ZN(I17898) );
INV_X32 U_g10995 ( .A(I17898), .ZN(g10995) );
INV_X32 U_I17901 ( .A(g6369), .ZN(I17901) );
INV_X32 U_g10996 ( .A(I17901), .ZN(g10996) );
INV_X32 U_I17904 ( .A(g6713), .ZN(I17904) );
INV_X32 U_g10999 ( .A(I17904), .ZN(g10999) );
INV_X32 U_I17907 ( .A(g5824), .ZN(I17907) );
INV_X32 U_g11002 ( .A(I17907), .ZN(g11002) );
INV_X32 U_I17910 ( .A(g7532), .ZN(I17910) );
INV_X32 U_g11003 ( .A(I17910), .ZN(g11003) );
INV_X32 U_I17913 ( .A(g7015), .ZN(I17913) );
INV_X32 U_g11004 ( .A(I17913), .ZN(g11004) );
INV_X32 U_I17916 ( .A(g7560), .ZN(I17916) );
INV_X32 U_g11007 ( .A(I17916), .ZN(g11007) );
INV_X32 U_I17919 ( .A(g7976), .ZN(I17919) );
INV_X32 U_g11008 ( .A(I17919), .ZN(g11008) );
INV_X32 U_I17922 ( .A(g8031), .ZN(I17922) );
INV_X32 U_g11011 ( .A(I17922), .ZN(g11011) );
INV_X32 U_I17925 ( .A(g7976), .ZN(I17925) );
INV_X32 U_g11014 ( .A(I17925), .ZN(g11014) );
INV_X32 U_I17928 ( .A(g8031), .ZN(I17928) );
INV_X32 U_g11017 ( .A(I17928), .ZN(g11017) );
INV_X32 U_g11020 ( .A(g6029), .ZN(g11020) );
INV_X32 U_g11021 ( .A(g6030), .ZN(g11021) );
INV_X32 U_I17933 ( .A(g3254), .ZN(I17933) );
INV_X32 U_g11022 ( .A(I17933), .ZN(g11022) );
INV_X32 U_I17936 ( .A(g6314), .ZN(I17936) );
INV_X32 U_g11025 ( .A(I17936), .ZN(g11025) );
INV_X32 U_I17939 ( .A(g6232), .ZN(I17939) );
INV_X32 U_g11028 ( .A(I17939), .ZN(g11028) );
INV_X32 U_I17942 ( .A(g5548), .ZN(I17942) );
INV_X32 U_g11031 ( .A(I17942), .ZN(g11031) );
INV_X32 U_I17945 ( .A(g5668), .ZN(I17945) );
INV_X32 U_g11032 ( .A(I17945), .ZN(g11032) );
INV_X32 U_I17948 ( .A(g6643), .ZN(I17948) );
INV_X32 U_g11035 ( .A(I17948), .ZN(g11035) );
INV_X32 U_I17951 ( .A(g6519), .ZN(I17951) );
INV_X32 U_g11036 ( .A(I17951), .ZN(g11036) );
INV_X32 U_I17954 ( .A(g6369), .ZN(I17954) );
INV_X32 U_g11039 ( .A(I17954), .ZN(g11039) );
INV_X32 U_I17957 ( .A(g6713), .ZN(I17957) );
INV_X32 U_g11042 ( .A(I17957), .ZN(g11042) );
INV_X32 U_I17960 ( .A(g6945), .ZN(I17960) );
INV_X32 U_g11045 ( .A(I17960), .ZN(g11045) );
INV_X32 U_I17963 ( .A(g6574), .ZN(I17963) );
INV_X32 U_g11048 ( .A(I17963), .ZN(g11048) );
INV_X32 U_I17966 ( .A(g7015), .ZN(I17966) );
INV_X32 U_g11051 ( .A(I17966), .ZN(g11051) );
INV_X32 U_I17969 ( .A(g5880), .ZN(I17969) );
INV_X32 U_g11054 ( .A(I17969), .ZN(g11054) );
INV_X32 U_I17972 ( .A(g7558), .ZN(I17972) );
INV_X32 U_g11055 ( .A(I17972), .ZN(g11055) );
INV_X32 U_I17975 ( .A(g7265), .ZN(I17975) );
INV_X32 U_g11056 ( .A(I17975), .ZN(g11056) );
INV_X32 U_I17978 ( .A(g7795), .ZN(I17978) );
INV_X32 U_g11059 ( .A(I17978), .ZN(g11059) );
INV_X32 U_I17981 ( .A(g7976), .ZN(I17981) );
INV_X32 U_g11063 ( .A(I17981), .ZN(g11063) );
INV_X32 U_I17984 ( .A(g7976), .ZN(I17984) );
INV_X32 U_g11066 ( .A(I17984), .ZN(g11066) );
INV_X32 U_g11069 ( .A(g8257), .ZN(g11069) );
INV_X32 U_g11078 ( .A(g6041), .ZN(g11078) );
INV_X32 U_I17989 ( .A(g3254), .ZN(I17989) );
INV_X32 U_g11079 ( .A(I17989), .ZN(g11079) );
INV_X32 U_I17992 ( .A(g6314), .ZN(I17992) );
INV_X32 U_g11082 ( .A(I17992), .ZN(g11082) );
INV_X32 U_I17995 ( .A(g6232), .ZN(I17995) );
INV_X32 U_g11085 ( .A(I17995), .ZN(g11085) );
INV_X32 U_I17998 ( .A(g5668), .ZN(I17998) );
INV_X32 U_g11088 ( .A(I17998), .ZN(g11088) );
INV_X32 U_I18001 ( .A(g6643), .ZN(I18001) );
INV_X32 U_g11091 ( .A(I18001), .ZN(g11091) );
INV_X32 U_I18004 ( .A(g3410), .ZN(I18004) );
INV_X32 U_g11092 ( .A(I18004), .ZN(g11092) );
INV_X32 U_I18007 ( .A(g6519), .ZN(I18007) );
INV_X32 U_g11095 ( .A(I18007), .ZN(g11095) );
INV_X32 U_I18010 ( .A(g6369), .ZN(I18010) );
INV_X32 U_g11098 ( .A(I18010), .ZN(g11098) );
INV_X32 U_I18013 ( .A(g5594), .ZN(I18013) );
INV_X32 U_g11101 ( .A(I18013), .ZN(g11101) );
INV_X32 U_I18016 ( .A(g5720), .ZN(I18016) );
INV_X32 U_g11102 ( .A(I18016), .ZN(g11102) );
INV_X32 U_I18019 ( .A(g6945), .ZN(I18019) );
INV_X32 U_g11105 ( .A(I18019), .ZN(g11105) );
INV_X32 U_I18022 ( .A(g6783), .ZN(I18022) );
INV_X32 U_g11108 ( .A(I18022), .ZN(g11108) );
INV_X32 U_I18025 ( .A(g6574), .ZN(I18025) );
INV_X32 U_g11111 ( .A(I18025), .ZN(g11111) );
INV_X32 U_I18028 ( .A(g7015), .ZN(I18028) );
INV_X32 U_g11114 ( .A(I18028), .ZN(g11114) );
INV_X32 U_I18031 ( .A(g7195), .ZN(I18031) );
INV_X32 U_g11117 ( .A(I18031), .ZN(g11117) );
INV_X32 U_I18034 ( .A(g6838), .ZN(I18034) );
INV_X32 U_g11120 ( .A(I18034), .ZN(g11120) );
INV_X32 U_I18037 ( .A(g7265), .ZN(I18037) );
INV_X32 U_g11123 ( .A(I18037), .ZN(g11123) );
INV_X32 U_I18040 ( .A(g7976), .ZN(I18040) );
INV_X32 U_g11126 ( .A(I18040), .ZN(g11126) );
INV_X32 U_I18043 ( .A(g7976), .ZN(I18043) );
INV_X32 U_g11129 ( .A(I18043), .ZN(g11129) );
INV_X32 U_I18046 ( .A(g3254), .ZN(I18046) );
INV_X32 U_g11132 ( .A(I18046), .ZN(g11132) );
INV_X32 U_I18049 ( .A(g6314), .ZN(I18049) );
INV_X32 U_g11135 ( .A(I18049), .ZN(g11135) );
INV_X32 U_I18052 ( .A(g6232), .ZN(I18052) );
INV_X32 U_g11138 ( .A(I18052), .ZN(g11138) );
INV_X32 U_I18055 ( .A(g5668), .ZN(I18055) );
INV_X32 U_g11141 ( .A(I18055), .ZN(g11141) );
INV_X32 U_I18058 ( .A(g6643), .ZN(I18058) );
INV_X32 U_g11144 ( .A(I18058), .ZN(g11144) );
INV_X32 U_I18061 ( .A(g3410), .ZN(I18061) );
INV_X32 U_g11145 ( .A(I18061), .ZN(g11145) );
INV_X32 U_I18064 ( .A(g6519), .ZN(I18064) );
INV_X32 U_g11148 ( .A(I18064), .ZN(g11148) );
INV_X32 U_I18067 ( .A(g6369), .ZN(I18067) );
INV_X32 U_g11151 ( .A(I18067), .ZN(g11151) );
INV_X32 U_I18070 ( .A(g5720), .ZN(I18070) );
INV_X32 U_g11154 ( .A(I18070), .ZN(g11154) );
INV_X32 U_I18073 ( .A(g6945), .ZN(I18073) );
INV_X32 U_g11157 ( .A(I18073), .ZN(g11157) );
INV_X32 U_I18076 ( .A(g3566), .ZN(I18076) );
INV_X32 U_g11160 ( .A(I18076), .ZN(g11160) );
INV_X32 U_I18079 ( .A(g6783), .ZN(I18079) );
INV_X32 U_g11163 ( .A(I18079), .ZN(g11163) );
INV_X32 U_I18082 ( .A(g6574), .ZN(I18082) );
INV_X32 U_g11166 ( .A(I18082), .ZN(g11166) );
INV_X32 U_I18085 ( .A(g5611), .ZN(I18085) );
INV_X32 U_g11169 ( .A(I18085), .ZN(g11169) );
INV_X32 U_I18088 ( .A(g5778), .ZN(I18088) );
INV_X32 U_g11170 ( .A(I18088), .ZN(g11170) );
INV_X32 U_I18091 ( .A(g7195), .ZN(I18091) );
INV_X32 U_g11173 ( .A(I18091), .ZN(g11173) );
INV_X32 U_I18094 ( .A(g7085), .ZN(I18094) );
INV_X32 U_g11176 ( .A(I18094), .ZN(g11176) );
INV_X32 U_I18097 ( .A(g6838), .ZN(I18097) );
INV_X32 U_g11179 ( .A(I18097), .ZN(g11179) );
INV_X32 U_I18100 ( .A(g7265), .ZN(I18100) );
INV_X32 U_g11182 ( .A(I18100), .ZN(g11182) );
INV_X32 U_I18103 ( .A(g7391), .ZN(I18103) );
INV_X32 U_g11185 ( .A(I18103), .ZN(g11185) );
INV_X32 U_g11190 ( .A(g3999), .ZN(g11190) );
INV_X32 U_I18121 ( .A(g3254), .ZN(I18121) );
INV_X32 U_g11199 ( .A(I18121), .ZN(g11199) );
INV_X32 U_I18124 ( .A(g6314), .ZN(I18124) );
INV_X32 U_g11202 ( .A(I18124), .ZN(g11202) );
INV_X32 U_I18127 ( .A(g6232), .ZN(I18127) );
INV_X32 U_g11205 ( .A(I18127), .ZN(g11205) );
INV_X32 U_I18130 ( .A(g5547), .ZN(I18130) );
INV_X32 U_g11208 ( .A(I18130), .ZN(g11208) );
INV_X32 U_I18133 ( .A(g6448), .ZN(I18133) );
INV_X32 U_g11209 ( .A(I18133), .ZN(g11209) );
INV_X32 U_I18136 ( .A(g5668), .ZN(I18136) );
INV_X32 U_g11210 ( .A(I18136), .ZN(g11210) );
INV_X32 U_I18139 ( .A(g6643), .ZN(I18139) );
INV_X32 U_g11213 ( .A(I18139), .ZN(g11213) );
INV_X32 U_I18142 ( .A(g3410), .ZN(I18142) );
INV_X32 U_g11216 ( .A(I18142), .ZN(g11216) );
INV_X32 U_I18145 ( .A(g6519), .ZN(I18145) );
INV_X32 U_g11219 ( .A(I18145), .ZN(g11219) );
INV_X32 U_I18148 ( .A(g6369), .ZN(I18148) );
INV_X32 U_g11222 ( .A(I18148), .ZN(g11222) );
INV_X32 U_I18151 ( .A(g5720), .ZN(I18151) );
INV_X32 U_g11225 ( .A(I18151), .ZN(g11225) );
INV_X32 U_I18154 ( .A(g6945), .ZN(I18154) );
INV_X32 U_g11228 ( .A(I18154), .ZN(g11228) );
INV_X32 U_I18157 ( .A(g3566), .ZN(I18157) );
INV_X32 U_g11231 ( .A(I18157), .ZN(g11231) );
INV_X32 U_I18160 ( .A(g6783), .ZN(I18160) );
INV_X32 U_g11234 ( .A(I18160), .ZN(g11234) );
INV_X32 U_I18163 ( .A(g6574), .ZN(I18163) );
INV_X32 U_g11237 ( .A(I18163), .ZN(g11237) );
INV_X32 U_I18166 ( .A(g5778), .ZN(I18166) );
INV_X32 U_g11240 ( .A(I18166), .ZN(g11240) );
INV_X32 U_I18169 ( .A(g7195), .ZN(I18169) );
INV_X32 U_g11243 ( .A(I18169), .ZN(g11243) );
INV_X32 U_I18172 ( .A(g3722), .ZN(I18172) );
INV_X32 U_g11246 ( .A(I18172), .ZN(g11246) );
INV_X32 U_I18175 ( .A(g7085), .ZN(I18175) );
INV_X32 U_g11249 ( .A(I18175), .ZN(g11249) );
INV_X32 U_I18178 ( .A(g6838), .ZN(I18178) );
INV_X32 U_g11252 ( .A(I18178), .ZN(g11252) );
INV_X32 U_I18181 ( .A(g5636), .ZN(I18181) );
INV_X32 U_g11255 ( .A(I18181), .ZN(g11255) );
INV_X32 U_I18184 ( .A(g5837), .ZN(I18184) );
INV_X32 U_g11256 ( .A(I18184), .ZN(g11256) );
INV_X32 U_I18187 ( .A(g7391), .ZN(I18187) );
INV_X32 U_g11259 ( .A(I18187), .ZN(g11259) );
INV_X32 U_I18211 ( .A(g6232), .ZN(I18211) );
INV_X32 U_g11265 ( .A(I18211), .ZN(g11265) );
INV_X32 U_I18214 ( .A(g3254), .ZN(I18214) );
INV_X32 U_g11268 ( .A(I18214), .ZN(g11268) );
INV_X32 U_I18217 ( .A(g6314), .ZN(I18217) );
INV_X32 U_g11271 ( .A(I18217), .ZN(g11271) );
INV_X32 U_I18220 ( .A(g6232), .ZN(I18220) );
INV_X32 U_g11274 ( .A(I18220), .ZN(g11274) );
INV_X32 U_I18223 ( .A(g6448), .ZN(I18223) );
INV_X32 U_g11277 ( .A(I18223), .ZN(g11277) );
INV_X32 U_I18226 ( .A(g5668), .ZN(I18226) );
INV_X32 U_g11278 ( .A(I18226), .ZN(g11278) );
INV_X32 U_I18229 ( .A(g3410), .ZN(I18229) );
INV_X32 U_g11281 ( .A(I18229), .ZN(g11281) );
INV_X32 U_I18232 ( .A(g6519), .ZN(I18232) );
INV_X32 U_g11284 ( .A(I18232), .ZN(g11284) );
INV_X32 U_I18235 ( .A(g6369), .ZN(I18235) );
INV_X32 U_g11287 ( .A(I18235), .ZN(g11287) );
INV_X32 U_I18238 ( .A(g5593), .ZN(I18238) );
INV_X32 U_g11290 ( .A(I18238), .ZN(g11290) );
INV_X32 U_I18241 ( .A(g6713), .ZN(I18241) );
INV_X32 U_g11291 ( .A(I18241), .ZN(g11291) );
INV_X32 U_I18244 ( .A(g5720), .ZN(I18244) );
INV_X32 U_g11294 ( .A(I18244), .ZN(g11294) );
INV_X32 U_I18247 ( .A(g6945), .ZN(I18247) );
INV_X32 U_g11297 ( .A(I18247), .ZN(g11297) );
INV_X32 U_I18250 ( .A(g3566), .ZN(I18250) );
INV_X32 U_g11300 ( .A(I18250), .ZN(g11300) );
INV_X32 U_I18253 ( .A(g6783), .ZN(I18253) );
INV_X32 U_g11303 ( .A(I18253), .ZN(g11303) );
INV_X32 U_I18256 ( .A(g6574), .ZN(I18256) );
INV_X32 U_g11306 ( .A(I18256), .ZN(g11306) );
INV_X32 U_I18259 ( .A(g5778), .ZN(I18259) );
INV_X32 U_g11309 ( .A(I18259), .ZN(g11309) );
INV_X32 U_I18262 ( .A(g7195), .ZN(I18262) );
INV_X32 U_g11312 ( .A(I18262), .ZN(g11312) );
INV_X32 U_I18265 ( .A(g3722), .ZN(I18265) );
INV_X32 U_g11315 ( .A(I18265), .ZN(g11315) );
INV_X32 U_I18268 ( .A(g7085), .ZN(I18268) );
INV_X32 U_g11318 ( .A(I18268), .ZN(g11318) );
INV_X32 U_I18271 ( .A(g6838), .ZN(I18271) );
INV_X32 U_g11321 ( .A(I18271), .ZN(g11321) );
INV_X32 U_I18274 ( .A(g5837), .ZN(I18274) );
INV_X32 U_g11324 ( .A(I18274), .ZN(g11324) );
INV_X32 U_I18277 ( .A(g7391), .ZN(I18277) );
INV_X32 U_g11327 ( .A(I18277), .ZN(g11327) );
INV_X32 U_g11332 ( .A(g4094), .ZN(g11332) );
INV_X32 U_I18295 ( .A(g6314), .ZN(I18295) );
INV_X32 U_g11341 ( .A(I18295), .ZN(g11341) );
INV_X32 U_I18298 ( .A(g6232), .ZN(I18298) );
INV_X32 U_g11344 ( .A(I18298), .ZN(g11344) );
INV_X32 U_I18302 ( .A(g3254), .ZN(I18302) );
INV_X32 U_g11348 ( .A(I18302), .ZN(g11348) );
INV_X32 U_I18305 ( .A(g6314), .ZN(I18305) );
INV_X32 U_g11351 ( .A(I18305), .ZN(g11351) );
INV_X32 U_I18308 ( .A(g6448), .ZN(I18308) );
INV_X32 U_g11354 ( .A(I18308), .ZN(g11354) );
INV_X32 U_I18311 ( .A(g5668), .ZN(I18311) );
INV_X32 U_g11355 ( .A(I18311), .ZN(g11355) );
INV_X32 U_I18314 ( .A(g6369), .ZN(I18314) );
INV_X32 U_g11358 ( .A(I18314), .ZN(g11358) );
INV_X32 U_I18317 ( .A(g3410), .ZN(I18317) );
INV_X32 U_g11361 ( .A(I18317), .ZN(g11361) );
INV_X32 U_I18320 ( .A(g6519), .ZN(I18320) );
INV_X32 U_g11364 ( .A(I18320), .ZN(g11364) );
INV_X32 U_I18323 ( .A(g6369), .ZN(I18323) );
INV_X32 U_g11367 ( .A(I18323), .ZN(g11367) );
INV_X32 U_I18326 ( .A(g6713), .ZN(I18326) );
INV_X32 U_g11370 ( .A(I18326), .ZN(g11370) );
INV_X32 U_I18329 ( .A(g5720), .ZN(I18329) );
INV_X32 U_g11373 ( .A(I18329), .ZN(g11373) );
INV_X32 U_I18332 ( .A(g3566), .ZN(I18332) );
INV_X32 U_g11376 ( .A(I18332), .ZN(g11376) );
INV_X32 U_I18335 ( .A(g6783), .ZN(I18335) );
INV_X32 U_g11379 ( .A(I18335), .ZN(g11379) );
INV_X32 U_I18338 ( .A(g6574), .ZN(I18338) );
INV_X32 U_g11382 ( .A(I18338), .ZN(g11382) );
INV_X32 U_I18341 ( .A(g5610), .ZN(I18341) );
INV_X32 U_g11385 ( .A(I18341), .ZN(g11385) );
INV_X32 U_I18344 ( .A(g7015), .ZN(I18344) );
INV_X32 U_g11386 ( .A(I18344), .ZN(g11386) );
INV_X32 U_I18347 ( .A(g5778), .ZN(I18347) );
INV_X32 U_g11389 ( .A(I18347), .ZN(g11389) );
INV_X32 U_I18350 ( .A(g7195), .ZN(I18350) );
INV_X32 U_g11392 ( .A(I18350), .ZN(g11392) );
INV_X32 U_I18353 ( .A(g3722), .ZN(I18353) );
INV_X32 U_g11395 ( .A(I18353), .ZN(g11395) );
INV_X32 U_I18356 ( .A(g7085), .ZN(I18356) );
INV_X32 U_g11398 ( .A(I18356), .ZN(g11398) );
INV_X32 U_I18359 ( .A(g6838), .ZN(I18359) );
INV_X32 U_g11401 ( .A(I18359), .ZN(g11401) );
INV_X32 U_I18362 ( .A(g5837), .ZN(I18362) );
INV_X32 U_g11404 ( .A(I18362), .ZN(g11404) );
INV_X32 U_I18365 ( .A(g7391), .ZN(I18365) );
INV_X32 U_g11407 ( .A(I18365), .ZN(g11407) );
INV_X32 U_I18375 ( .A(g3254), .ZN(I18375) );
INV_X32 U_g11411 ( .A(I18375), .ZN(g11411) );
INV_X32 U_I18378 ( .A(g6314), .ZN(I18378) );
INV_X32 U_g11414 ( .A(I18378), .ZN(g11414) );
INV_X32 U_I18381 ( .A(g6232), .ZN(I18381) );
INV_X32 U_g11417 ( .A(I18381), .ZN(g11417) );
INV_X32 U_I18386 ( .A(g3254), .ZN(I18386) );
INV_X32 U_g11422 ( .A(I18386), .ZN(g11422) );
INV_X32 U_I18389 ( .A(g6519), .ZN(I18389) );
INV_X32 U_g11425 ( .A(I18389), .ZN(g11425) );
INV_X32 U_I18392 ( .A(g6369), .ZN(I18392) );
INV_X32 U_g11428 ( .A(I18392), .ZN(g11428) );
INV_X32 U_I18396 ( .A(g3410), .ZN(I18396) );
INV_X32 U_g11432 ( .A(I18396), .ZN(g11432) );
INV_X32 U_I18399 ( .A(g6519), .ZN(I18399) );
INV_X32 U_g11435 ( .A(I18399), .ZN(g11435) );
INV_X32 U_I18402 ( .A(g6713), .ZN(I18402) );
INV_X32 U_g11438 ( .A(I18402), .ZN(g11438) );
INV_X32 U_I18405 ( .A(g5720), .ZN(I18405) );
INV_X32 U_g11441 ( .A(I18405), .ZN(g11441) );
INV_X32 U_I18408 ( .A(g6574), .ZN(I18408) );
INV_X32 U_g11444 ( .A(I18408), .ZN(g11444) );
INV_X32 U_I18411 ( .A(g3566), .ZN(I18411) );
INV_X32 U_g11447 ( .A(I18411), .ZN(g11447) );
INV_X32 U_I18414 ( .A(g6783), .ZN(I18414) );
INV_X32 U_g11450 ( .A(I18414), .ZN(g11450) );
INV_X32 U_I18417 ( .A(g6574), .ZN(I18417) );
INV_X32 U_g11453 ( .A(I18417), .ZN(g11453) );
INV_X32 U_I18420 ( .A(g7015), .ZN(I18420) );
INV_X32 U_g11456 ( .A(I18420), .ZN(g11456) );
INV_X32 U_I18423 ( .A(g5778), .ZN(I18423) );
INV_X32 U_g11459 ( .A(I18423), .ZN(g11459) );
INV_X32 U_I18426 ( .A(g3722), .ZN(I18426) );
INV_X32 U_g11462 ( .A(I18426), .ZN(g11462) );
INV_X32 U_I18429 ( .A(g7085), .ZN(I18429) );
INV_X32 U_g11465 ( .A(I18429), .ZN(g11465) );
INV_X32 U_I18432 ( .A(g6838), .ZN(I18432) );
INV_X32 U_g11468 ( .A(I18432), .ZN(g11468) );
INV_X32 U_I18435 ( .A(g5635), .ZN(I18435) );
INV_X32 U_g11471 ( .A(I18435), .ZN(g11471) );
INV_X32 U_I18438 ( .A(g7265), .ZN(I18438) );
INV_X32 U_g11472 ( .A(I18438), .ZN(g11472) );
INV_X32 U_I18441 ( .A(g5837), .ZN(I18441) );
INV_X32 U_g11475 ( .A(I18441), .ZN(g11475) );
INV_X32 U_I18444 ( .A(g7391), .ZN(I18444) );
INV_X32 U_g11478 ( .A(I18444), .ZN(g11478) );
INV_X32 U_g11481 ( .A(g4204), .ZN(g11481) );
INV_X32 U_g11490 ( .A(g8276), .ZN(g11490) );
INV_X32 U_I18449 ( .A(g10868), .ZN(I18449) );
INV_X32 U_g11491 ( .A(I18449), .ZN(g11491) );
INV_X32 U_I18452 ( .A(g10930), .ZN(I18452) );
INV_X32 U_g11492 ( .A(I18452), .ZN(g11492) );
INV_X32 U_I18455 ( .A(g11031), .ZN(I18455) );
INV_X32 U_g11493 ( .A(I18455), .ZN(g11493) );
INV_X32 U_I18458 ( .A(g11208), .ZN(I18458) );
INV_X32 U_g11494 ( .A(I18458), .ZN(g11494) );
INV_X32 U_I18461 ( .A(g10931), .ZN(I18461) );
INV_X32 U_g11495 ( .A(I18461), .ZN(g11495) );
INV_X32 U_I18464 ( .A(g8620), .ZN(I18464) );
INV_X32 U_g11496 ( .A(I18464), .ZN(g11496) );
INV_X32 U_I18467 ( .A(g8769), .ZN(I18467) );
INV_X32 U_g11497 ( .A(I18467), .ZN(g11497) );
INV_X32 U_I18470 ( .A(g8808), .ZN(I18470) );
INV_X32 U_g11498 ( .A(I18470), .ZN(g11498) );
INV_X32 U_I18473 ( .A(g8839), .ZN(I18473) );
INV_X32 U_g11499 ( .A(I18473), .ZN(g11499) );
INV_X32 U_I18476 ( .A(g8791), .ZN(I18476) );
INV_X32 U_g11500 ( .A(I18476), .ZN(g11500) );
INV_X32 U_I18479 ( .A(g8820), .ZN(I18479) );
INV_X32 U_g11501 ( .A(I18479), .ZN(g11501) );
INV_X32 U_I18482 ( .A(g8859), .ZN(I18482) );
INV_X32 U_g11502 ( .A(I18482), .ZN(g11502) );
INV_X32 U_I18485 ( .A(g8809), .ZN(I18485) );
INV_X32 U_g11503 ( .A(I18485), .ZN(g11503) );
INV_X32 U_I18488 ( .A(g8840), .ZN(I18488) );
INV_X32 U_g11504 ( .A(I18488), .ZN(g11504) );
INV_X32 U_I18491 ( .A(g8891), .ZN(I18491) );
INV_X32 U_g11505 ( .A(I18491), .ZN(g11505) );
INV_X32 U_I18494 ( .A(g8821), .ZN(I18494) );
INV_X32 U_g11506 ( .A(I18494), .ZN(g11506) );
INV_X32 U_I18497 ( .A(g8860), .ZN(I18497) );
INV_X32 U_g11507 ( .A(I18497), .ZN(g11507) );
INV_X32 U_I18500 ( .A(g8924), .ZN(I18500) );
INV_X32 U_g11508 ( .A(I18500), .ZN(g11508) );
INV_X32 U_I18503 ( .A(g8658), .ZN(I18503) );
INV_X32 U_g11509 ( .A(I18503), .ZN(g11509) );
INV_X32 U_I18506 ( .A(g8699), .ZN(I18506) );
INV_X32 U_g11510 ( .A(I18506), .ZN(g11510) );
INV_X32 U_I18509 ( .A(g8770), .ZN(I18509) );
INV_X32 U_g11511 ( .A(I18509), .ZN(g11511) );
INV_X32 U_I18512 ( .A(g9309), .ZN(I18512) );
INV_X32 U_g11512 ( .A(I18512), .ZN(g11512) );
INV_X32 U_I18515 ( .A(g8843), .ZN(I18515) );
INV_X32 U_g11513 ( .A(I18515), .ZN(g11513) );
INV_X32 U_I18518 ( .A(g8893), .ZN(I18518) );
INV_X32 U_g11514 ( .A(I18518), .ZN(g11514) );
INV_X32 U_I18521 ( .A(g9449), .ZN(I18521) );
INV_X32 U_g11515 ( .A(I18521), .ZN(g11515) );
INV_X32 U_I18524 ( .A(g9640), .ZN(I18524) );
INV_X32 U_g11516 ( .A(I18524), .ZN(g11516) );
INV_X32 U_I18527 ( .A(g10017), .ZN(I18527) );
INV_X32 U_g11517 ( .A(I18527), .ZN(g11517) );
INV_X32 U_I18530 ( .A(g10888), .ZN(I18530) );
INV_X32 U_g11518 ( .A(I18530), .ZN(g11518) );
INV_X32 U_I18533 ( .A(g10967), .ZN(I18533) );
INV_X32 U_g11519 ( .A(I18533), .ZN(g11519) );
INV_X32 U_I18536 ( .A(g11101), .ZN(I18536) );
INV_X32 U_g11520 ( .A(I18536), .ZN(g11520) );
INV_X32 U_I18539 ( .A(g11290), .ZN(I18539) );
INV_X32 U_g11521 ( .A(I18539), .ZN(g11521) );
INV_X32 U_I18542 ( .A(g10968), .ZN(I18542) );
INV_X32 U_g11522 ( .A(I18542), .ZN(g11522) );
INV_X32 U_I18545 ( .A(g8630), .ZN(I18545) );
INV_X32 U_g11523 ( .A(I18545), .ZN(g11523) );
INV_X32 U_I18548 ( .A(g8792), .ZN(I18548) );
INV_X32 U_g11524 ( .A(I18548), .ZN(g11524) );
INV_X32 U_I18551 ( .A(g8824), .ZN(I18551) );
INV_X32 U_g11525 ( .A(I18551), .ZN(g11525) );
INV_X32 U_I18554 ( .A(g8866), .ZN(I18554) );
INV_X32 U_g11526 ( .A(I18554), .ZN(g11526) );
INV_X32 U_I18557 ( .A(g8810), .ZN(I18557) );
INV_X32 U_g11527 ( .A(I18557), .ZN(g11527) );
INV_X32 U_I18560 ( .A(g8844), .ZN(I18560) );
INV_X32 U_g11528 ( .A(I18560), .ZN(g11528) );
INV_X32 U_I18563 ( .A(g8897), .ZN(I18563) );
INV_X32 U_g11529 ( .A(I18563), .ZN(g11529) );
INV_X32 U_I18566 ( .A(g8825), .ZN(I18566) );
INV_X32 U_g11530 ( .A(I18566), .ZN(g11530) );
INV_X32 U_I18569 ( .A(g8867), .ZN(I18569) );
INV_X32 U_g11531 ( .A(I18569), .ZN(g11531) );
INV_X32 U_I18572 ( .A(g8931), .ZN(I18572) );
INV_X32 U_g11532 ( .A(I18572), .ZN(g11532) );
INV_X32 U_I18575 ( .A(g8845), .ZN(I18575) );
INV_X32 U_g11533 ( .A(I18575), .ZN(g11533) );
INV_X32 U_I18578 ( .A(g8898), .ZN(I18578) );
INV_X32 U_g11534 ( .A(I18578), .ZN(g11534) );
INV_X32 U_I18581 ( .A(g8964), .ZN(I18581) );
INV_X32 U_g11535 ( .A(I18581), .ZN(g11535) );
INV_X32 U_I18584 ( .A(g8677), .ZN(I18584) );
INV_X32 U_g11536 ( .A(I18584), .ZN(g11536) );
INV_X32 U_I18587 ( .A(g8718), .ZN(I18587) );
INV_X32 U_g11537 ( .A(I18587), .ZN(g11537) );
INV_X32 U_I18590 ( .A(g8793), .ZN(I18590) );
INV_X32 U_g11538 ( .A(I18590), .ZN(g11538) );
INV_X32 U_I18593 ( .A(g9390), .ZN(I18593) );
INV_X32 U_g11539 ( .A(I18593), .ZN(g11539) );
INV_X32 U_I18596 ( .A(g8870), .ZN(I18596) );
INV_X32 U_g11540 ( .A(I18596), .ZN(g11540) );
INV_X32 U_I18599 ( .A(g8933), .ZN(I18599) );
INV_X32 U_g11541 ( .A(I18599), .ZN(g11541) );
INV_X32 U_I18602 ( .A(g9591), .ZN(I18602) );
INV_X32 U_g11542 ( .A(I18602), .ZN(g11542) );
INV_X32 U_I18605 ( .A(g9786), .ZN(I18605) );
INV_X32 U_g11543 ( .A(I18605), .ZN(g11543) );
INV_X32 U_I18608 ( .A(g10126), .ZN(I18608) );
INV_X32 U_g11544 ( .A(I18608), .ZN(g11544) );
INV_X32 U_I18611 ( .A(g10909), .ZN(I18611) );
INV_X32 U_g11545 ( .A(I18611), .ZN(g11545) );
INV_X32 U_I18614 ( .A(g11002), .ZN(I18614) );
INV_X32 U_g11546 ( .A(I18614), .ZN(g11546) );
INV_X32 U_I18617 ( .A(g11169), .ZN(I18617) );
INV_X32 U_g11547 ( .A(I18617), .ZN(g11547) );
INV_X32 U_I18620 ( .A(g11385), .ZN(I18620) );
INV_X32 U_g11548 ( .A(I18620), .ZN(g11548) );
INV_X32 U_I18623 ( .A(g11003), .ZN(I18623) );
INV_X32 U_g11549 ( .A(I18623), .ZN(g11549) );
INV_X32 U_I18626 ( .A(g8649), .ZN(I18626) );
INV_X32 U_g11550 ( .A(I18626), .ZN(g11550) );
INV_X32 U_I18629 ( .A(g8811), .ZN(I18629) );
INV_X32 U_g11551 ( .A(I18629), .ZN(g11551) );
INV_X32 U_I18632 ( .A(g8850), .ZN(I18632) );
INV_X32 U_g11552 ( .A(I18632), .ZN(g11552) );
INV_X32 U_I18635 ( .A(g8904), .ZN(I18635) );
INV_X32 U_g11553 ( .A(I18635), .ZN(g11553) );
INV_X32 U_I18638 ( .A(g8826), .ZN(I18638) );
INV_X32 U_g11554 ( .A(I18638), .ZN(g11554) );
INV_X32 U_I18641 ( .A(g8871), .ZN(I18641) );
INV_X32 U_g11555 ( .A(I18641), .ZN(g11555) );
INV_X32 U_I18644 ( .A(g8937), .ZN(I18644) );
INV_X32 U_g11556 ( .A(I18644), .ZN(g11556) );
INV_X32 U_I18647 ( .A(g8851), .ZN(I18647) );
INV_X32 U_g11557 ( .A(I18647), .ZN(g11557) );
INV_X32 U_I18650 ( .A(g8905), .ZN(I18650) );
INV_X32 U_g11558 ( .A(I18650), .ZN(g11558) );
INV_X32 U_I18653 ( .A(g8971), .ZN(I18653) );
INV_X32 U_g11559 ( .A(I18653), .ZN(g11559) );
INV_X32 U_I18656 ( .A(g8872), .ZN(I18656) );
INV_X32 U_g11560 ( .A(I18656), .ZN(g11560) );
INV_X32 U_I18659 ( .A(g8938), .ZN(I18659) );
INV_X32 U_g11561 ( .A(I18659), .ZN(g11561) );
INV_X32 U_I18662 ( .A(g8996), .ZN(I18662) );
INV_X32 U_g11562 ( .A(I18662), .ZN(g11562) );
INV_X32 U_I18665 ( .A(g8689), .ZN(I18665) );
INV_X32 U_g11563 ( .A(I18665), .ZN(g11563) );
INV_X32 U_I18668 ( .A(g8756), .ZN(I18668) );
INV_X32 U_g11564 ( .A(I18668), .ZN(g11564) );
INV_X32 U_I18671 ( .A(g8812), .ZN(I18671) );
INV_X32 U_g11565 ( .A(I18671), .ZN(g11565) );
INV_X32 U_I18674 ( .A(g9487), .ZN(I18674) );
INV_X32 U_g11566 ( .A(I18674), .ZN(g11566) );
INV_X32 U_I18677 ( .A(g8908), .ZN(I18677) );
INV_X32 U_g11567 ( .A(I18677), .ZN(g11567) );
INV_X32 U_I18680 ( .A(g8973), .ZN(I18680) );
INV_X32 U_g11568 ( .A(I18680), .ZN(g11568) );
INV_X32 U_I18683 ( .A(g9733), .ZN(I18683) );
INV_X32 U_g11569 ( .A(I18683), .ZN(g11569) );
INV_X32 U_I18686 ( .A(g9932), .ZN(I18686) );
INV_X32 U_g11570 ( .A(I18686), .ZN(g11570) );
INV_X32 U_I18689 ( .A(g10231), .ZN(I18689) );
INV_X32 U_g11571 ( .A(I18689), .ZN(g11571) );
INV_X32 U_I18692 ( .A(g10935), .ZN(I18692) );
INV_X32 U_g11572 ( .A(I18692), .ZN(g11572) );
INV_X32 U_I18695 ( .A(g11054), .ZN(I18695) );
INV_X32 U_g11573 ( .A(I18695), .ZN(g11573) );
INV_X32 U_I18698 ( .A(g11255), .ZN(I18698) );
INV_X32 U_g11574 ( .A(I18698), .ZN(g11574) );
INV_X32 U_I18701 ( .A(g11471), .ZN(I18701) );
INV_X32 U_g11575 ( .A(I18701), .ZN(g11575) );
INV_X32 U_I18704 ( .A(g11055), .ZN(I18704) );
INV_X32 U_g11576 ( .A(I18704), .ZN(g11576) );
INV_X32 U_I18707 ( .A(g8665), .ZN(I18707) );
INV_X32 U_g11577 ( .A(I18707), .ZN(g11577) );
INV_X32 U_I18710 ( .A(g8827), .ZN(I18710) );
INV_X32 U_g11578 ( .A(I18710), .ZN(g11578) );
INV_X32 U_I18713 ( .A(g8877), .ZN(I18713) );
INV_X32 U_g11579 ( .A(I18713), .ZN(g11579) );
INV_X32 U_I18716 ( .A(g8944), .ZN(I18716) );
INV_X32 U_g11580 ( .A(I18716), .ZN(g11580) );
INV_X32 U_I18719 ( .A(g8852), .ZN(I18719) );
INV_X32 U_g11581 ( .A(I18719), .ZN(g11581) );
INV_X32 U_I18722 ( .A(g8909), .ZN(I18722) );
INV_X32 U_g11582 ( .A(I18722), .ZN(g11582) );
INV_X32 U_I18725 ( .A(g8977), .ZN(I18725) );
INV_X32 U_g11583 ( .A(I18725), .ZN(g11583) );
INV_X32 U_I18728 ( .A(g8878), .ZN(I18728) );
INV_X32 U_g11584 ( .A(I18728), .ZN(g11584) );
INV_X32 U_I18731 ( .A(g8945), .ZN(I18731) );
INV_X32 U_g11585 ( .A(I18731), .ZN(g11585) );
INV_X32 U_I18734 ( .A(g9003), .ZN(I18734) );
INV_X32 U_g11586 ( .A(I18734), .ZN(g11586) );
INV_X32 U_I18737 ( .A(g8910), .ZN(I18737) );
INV_X32 U_g11587 ( .A(I18737), .ZN(g11587) );
INV_X32 U_I18740 ( .A(g8978), .ZN(I18740) );
INV_X32 U_g11588 ( .A(I18740), .ZN(g11588) );
INV_X32 U_I18743 ( .A(g9025), .ZN(I18743) );
INV_X32 U_g11589 ( .A(I18743), .ZN(g11589) );
INV_X32 U_I18746 ( .A(g8707), .ZN(I18746) );
INV_X32 U_g11590 ( .A(I18746), .ZN(g11590) );
INV_X32 U_I18749 ( .A(g8779), .ZN(I18749) );
INV_X32 U_g11591 ( .A(I18749), .ZN(g11591) );
INV_X32 U_I18752 ( .A(g8828), .ZN(I18752) );
INV_X32 U_g11592 ( .A(I18752), .ZN(g11592) );
INV_X32 U_I18755 ( .A(g9629), .ZN(I18755) );
INV_X32 U_g11593 ( .A(I18755), .ZN(g11593) );
INV_X32 U_I18758 ( .A(g8948), .ZN(I18758) );
INV_X32 U_g11594 ( .A(I18758), .ZN(g11594) );
INV_X32 U_I18761 ( .A(g9005), .ZN(I18761) );
INV_X32 U_g11595 ( .A(I18761), .ZN(g11595) );
INV_X32 U_I18764 ( .A(g9879), .ZN(I18764) );
INV_X32 U_g11596 ( .A(I18764), .ZN(g11596) );
INV_X32 U_I18767 ( .A(g10086), .ZN(I18767) );
INV_X32 U_g11597 ( .A(I18767), .ZN(g11597) );
INV_X32 U_I18770 ( .A(g10333), .ZN(I18770) );
INV_X32 U_g11598 ( .A(I18770), .ZN(g11598) );
INV_X32 U_I18773 ( .A(g10830), .ZN(I18773) );
INV_X32 U_g11599 ( .A(I18773), .ZN(g11599) );
INV_X32 U_I18777 ( .A(g9050), .ZN(I18777) );
INV_X32 U_g11603 ( .A(I18777), .ZN(g11603) );
INV_X32 U_I18780 ( .A(g10870), .ZN(I18780) );
INV_X32 U_g11606 ( .A(I18780), .ZN(g11606) );
INV_X32 U_I18784 ( .A(g9067), .ZN(I18784) );
INV_X32 U_g11608 ( .A(I18784), .ZN(g11608) );
INV_X32 U_I18787 ( .A(g10910), .ZN(I18787) );
INV_X32 U_g11611 ( .A(I18787), .ZN(g11611) );
INV_X32 U_I18791 ( .A(g9084), .ZN(I18791) );
INV_X32 U_g11613 ( .A(I18791), .ZN(g11613) );
INV_X32 U_I18794 ( .A(g10973), .ZN(I18794) );
INV_X32 U_g11616 ( .A(I18794), .ZN(g11616) );
INV_X32 U_g11620 ( .A(g10601), .ZN(g11620) );
INV_X32 U_g11623 ( .A(g10961), .ZN(g11623) );
INV_X32 U_I18810 ( .A(g10813), .ZN(I18810) );
INV_X32 U_g11628 ( .A(I18810), .ZN(g11628) );
INV_X32 U_I18813 ( .A(g10850), .ZN(I18813) );
INV_X32 U_g11629 ( .A(I18813), .ZN(g11629) );
INV_X32 U_I18817 ( .A(g9067), .ZN(I18817) );
INV_X32 U_g11633 ( .A(I18817), .ZN(g11633) );
INV_X32 U_I18820 ( .A(g10890), .ZN(I18820) );
INV_X32 U_g11636 ( .A(I18820), .ZN(g11636) );
INV_X32 U_I18824 ( .A(g9084), .ZN(I18824) );
INV_X32 U_g11638 ( .A(I18824), .ZN(g11638) );
INV_X32 U_I18827 ( .A(g10936), .ZN(I18827) );
INV_X32 U_g11641 ( .A(I18827), .ZN(g11641) );
INV_X32 U_g11642 ( .A(g10646), .ZN(g11642) );
INV_X32 U_I18835 ( .A(g10834), .ZN(I18835) );
INV_X32 U_g11651 ( .A(I18835), .ZN(g11651) );
INV_X32 U_I18838 ( .A(g10871), .ZN(I18838) );
INV_X32 U_g11652 ( .A(I18838), .ZN(g11652) );
INV_X32 U_I18842 ( .A(g9084), .ZN(I18842) );
INV_X32 U_g11656 ( .A(I18842), .ZN(g11656) );
INV_X32 U_I18845 ( .A(g10911), .ZN(I18845) );
INV_X32 U_g11659 ( .A(I18845), .ZN(g11659) );
INV_X32 U_I18854 ( .A(g10854), .ZN(I18854) );
INV_X32 U_g11670 ( .A(I18854), .ZN(g11670) );
INV_X32 U_I18857 ( .A(g10891), .ZN(I18857) );
INV_X32 U_g11671 ( .A(I18857), .ZN(g11671) );
INV_X32 U_I18866 ( .A(g10875), .ZN(I18866) );
INV_X32 U_g11682 ( .A(I18866), .ZN(g11682) );
INV_X32 U_g11706 ( .A(g10928), .ZN(g11706) );
INV_X32 U_g11732 ( .A(g10826), .ZN(g11732) );
INV_X32 U_g11734 ( .A(g10843), .ZN(g11734) );
INV_X32 U_g11735 ( .A(g10859), .ZN(g11735) );
INV_X32 U_g11736 ( .A(g10862), .ZN(g11736) );
INV_X32 U_g11737 ( .A(g10809), .ZN(g11737) );
INV_X32 U_g11740 ( .A(g10877), .ZN(g11740) );
INV_X32 U_g11741 ( .A(g10880), .ZN(g11741) );
INV_X32 U_g11742 ( .A(g10883), .ZN(g11742) );
INV_X32 U_g11743 ( .A(g8530), .ZN(g11743) );
INV_X32 U_g11745 ( .A(g10892), .ZN(g11745) );
INV_X32 U_g11746 ( .A(g10895), .ZN(g11746) );
INV_X32 U_g11747 ( .A(g10898), .ZN(g11747) );
INV_X32 U_g11748 ( .A(g10901), .ZN(g11748) );
INV_X32 U_I18929 ( .A(g10711), .ZN(I18929) );
INV_X32 U_g11749 ( .A(I18929), .ZN(g11749) );
INV_X32 U_g11758 ( .A(g8514), .ZN(g11758) );
INV_X32 U_g11761 ( .A(g10912), .ZN(g11761) );
INV_X32 U_g11762 ( .A(g10915), .ZN(g11762) );
INV_X32 U_g11763 ( .A(g10918), .ZN(g11763) );
INV_X32 U_g11764 ( .A(g10921), .ZN(g11764) );
INV_X32 U_g11765 ( .A(g10924), .ZN(g11765) );
INV_X32 U_g11766 ( .A(g10886), .ZN(g11766) );
INV_X32 U_I18943 ( .A(g9149), .ZN(I18943) );
INV_X32 U_g11769 ( .A(I18943), .ZN(g11769) );
INV_X32 U_g11770 ( .A(g10932), .ZN(g11770) );
INV_X32 U_g11774 ( .A(g10937), .ZN(g11774) );
INV_X32 U_g11775 ( .A(g10940), .ZN(g11775) );
INV_X32 U_g11776 ( .A(g10943), .ZN(g11776) );
INV_X32 U_g11777 ( .A(g10946), .ZN(g11777) );
INV_X32 U_g11778 ( .A(g10949), .ZN(g11778) );
INV_X32 U_g11779 ( .A(g10906), .ZN(g11779) );
INV_X32 U_g11782 ( .A(g10963), .ZN(g11782) );
INV_X32 U_g11783 ( .A(g10966), .ZN(g11783) );
INV_X32 U_I18962 ( .A(g9159), .ZN(I18962) );
INV_X32 U_g11786 ( .A(I18962), .ZN(g11786) );
INV_X32 U_g11787 ( .A(g10969), .ZN(g11787) );
INV_X32 U_I18969 ( .A(g8726), .ZN(I18969) );
INV_X32 U_g11791 ( .A(I18969), .ZN(g11791) );
INV_X32 U_g11794 ( .A(g10974), .ZN(g11794) );
INV_X32 U_g11795 ( .A(g10977), .ZN(g11795) );
INV_X32 U_g11796 ( .A(g10980), .ZN(g11796) );
INV_X32 U_g11797 ( .A(g10983), .ZN(g11797) );
INV_X32 U_g11798 ( .A(g10867), .ZN(g11798) );
INV_X32 U_g11801 ( .A(g10988), .ZN(g11801) );
INV_X32 U_g11802 ( .A(g10991), .ZN(g11802) );
INV_X32 U_g11803 ( .A(g10994), .ZN(g11803) );
INV_X32 U_g11804 ( .A(g10995), .ZN(g11804) );
INV_X32 U_g11808 ( .A(g10996), .ZN(g11808) );
INV_X32 U_g11809 ( .A(g10999), .ZN(g11809) );
INV_X32 U_I18990 ( .A(g9183), .ZN(I18990) );
INV_X32 U_g11812 ( .A(I18990), .ZN(g11812) );
INV_X32 U_g11813 ( .A(g11004), .ZN(g11813) );
INV_X32 U_g11817 ( .A(g11008), .ZN(g11817) );
INV_X32 U_g11818 ( .A(g11011), .ZN(g11818) );
INV_X32 U_g11819 ( .A(g11014), .ZN(g11819) );
INV_X32 U_g11820 ( .A(g11017), .ZN(g11820) );
INV_X32 U_g11821 ( .A(g10848), .ZN(g11821) );
INV_X32 U_g11824 ( .A(g11022), .ZN(g11824) );
INV_X32 U_g11825 ( .A(g11025), .ZN(g11825) );
INV_X32 U_g11826 ( .A(g11028), .ZN(g11826) );
INV_X32 U_g11827 ( .A(g11032), .ZN(g11827) );
INV_X32 U_g11829 ( .A(g11035), .ZN(g11829) );
INV_X32 U_g11834 ( .A(g11036), .ZN(g11834) );
INV_X32 U_g11835 ( .A(g11039), .ZN(g11835) );
INV_X32 U_g11836 ( .A(g11042), .ZN(g11836) );
INV_X32 U_g11837 ( .A(g11045), .ZN(g11837) );
INV_X32 U_g11841 ( .A(g11048), .ZN(g11841) );
INV_X32 U_g11842 ( .A(g11051), .ZN(g11842) );
INV_X32 U_I19025 ( .A(g9225), .ZN(I19025) );
INV_X32 U_g11845 ( .A(I19025), .ZN(g11845) );
INV_X32 U_g11846 ( .A(g11056), .ZN(g11846) );
INV_X32 U_I19030 ( .A(g8726), .ZN(I19030) );
INV_X32 U_g11848 ( .A(I19030), .ZN(g11848) );
INV_X32 U_g11852 ( .A(g11063), .ZN(g11852) );
INV_X32 U_g11853 ( .A(g11066), .ZN(g11853) );
INV_X32 U_g11854 ( .A(g11078), .ZN(g11854) );
INV_X32 U_g11856 ( .A(g11079), .ZN(g11856) );
INV_X32 U_g11857 ( .A(g11082), .ZN(g11857) );
INV_X32 U_g11858 ( .A(g11085), .ZN(g11858) );
INV_X32 U_g11859 ( .A(g11088), .ZN(g11859) );
INV_X32 U_g11862 ( .A(g11091), .ZN(g11862) );
INV_X32 U_g11866 ( .A(g11092), .ZN(g11866) );
INV_X32 U_g11867 ( .A(g11095), .ZN(g11867) );
INV_X32 U_g11868 ( .A(g11098), .ZN(g11868) );
INV_X32 U_g11869 ( .A(g11102), .ZN(g11869) );
INV_X32 U_g11871 ( .A(g11105), .ZN(g11871) );
INV_X32 U_g11876 ( .A(g11108), .ZN(g11876) );
INV_X32 U_g11877 ( .A(g11111), .ZN(g11877) );
INV_X32 U_g11878 ( .A(g11114), .ZN(g11878) );
INV_X32 U_g11879 ( .A(g11117), .ZN(g11879) );
INV_X32 U_g11883 ( .A(g11120), .ZN(g11883) );
INV_X32 U_g11884 ( .A(g11123), .ZN(g11884) );
INV_X32 U_g11886 ( .A(g11126), .ZN(g11886) );
INV_X32 U_g11887 ( .A(g11129), .ZN(g11887) );
INV_X32 U_g11888 ( .A(g11021), .ZN(g11888) );
INV_X32 U_g11891 ( .A(g11132), .ZN(g11891) );
INV_X32 U_g11892 ( .A(g11135), .ZN(g11892) );
INV_X32 U_g11893 ( .A(g11138), .ZN(g11893) );
INV_X32 U_g11894 ( .A(g11141), .ZN(g11894) );
INV_X32 U_g11895 ( .A(g11144), .ZN(g11895) );
INV_X32 U_g11898 ( .A(g11145), .ZN(g11898) );
INV_X32 U_g11899 ( .A(g11148), .ZN(g11899) );
INV_X32 U_g11900 ( .A(g11151), .ZN(g11900) );
INV_X32 U_g11901 ( .A(g11154), .ZN(g11901) );
INV_X32 U_g11904 ( .A(g11157), .ZN(g11904) );
INV_X32 U_g11908 ( .A(g11160), .ZN(g11908) );
INV_X32 U_g11909 ( .A(g11163), .ZN(g11909) );
INV_X32 U_g11910 ( .A(g11166), .ZN(g11910) );
INV_X32 U_g11911 ( .A(g11170), .ZN(g11911) );
INV_X32 U_g11913 ( .A(g11173), .ZN(g11913) );
INV_X32 U_g11918 ( .A(g11176), .ZN(g11918) );
INV_X32 U_g11919 ( .A(g11179), .ZN(g11919) );
INV_X32 U_g11920 ( .A(g11182), .ZN(g11920) );
INV_X32 U_g11921 ( .A(g11185), .ZN(g11921) );
INV_X32 U_I19105 ( .A(g8726), .ZN(I19105) );
INV_X32 U_g11923 ( .A(I19105), .ZN(g11923) );
INV_X32 U_g11927 ( .A(g10987), .ZN(g11927) );
INV_X32 U_g11929 ( .A(g11199), .ZN(g11929) );
INV_X32 U_g11930 ( .A(g11202), .ZN(g11930) );
INV_X32 U_g11931 ( .A(g11205), .ZN(g11931) );
INV_X32 U_g11932 ( .A(g11209), .ZN(g11932) );
INV_X32 U_g11933 ( .A(g11210), .ZN(g11933) );
INV_X32 U_g11936 ( .A(g11213), .ZN(g11936) );
INV_X32 U_I19119 ( .A(g9202), .ZN(I19119) );
INV_X32 U_g11937 ( .A(I19119), .ZN(g11937) );
INV_X32 U_g11941 ( .A(g11216), .ZN(g11941) );
INV_X32 U_g11942 ( .A(g11219), .ZN(g11942) );
INV_X32 U_g11943 ( .A(g11222), .ZN(g11943) );
INV_X32 U_g11944 ( .A(g11225), .ZN(g11944) );
INV_X32 U_g11945 ( .A(g11228), .ZN(g11945) );
INV_X32 U_g11948 ( .A(g11231), .ZN(g11948) );
INV_X32 U_g11949 ( .A(g11234), .ZN(g11949) );
INV_X32 U_g11950 ( .A(g11237), .ZN(g11950) );
INV_X32 U_g11951 ( .A(g11240), .ZN(g11951) );
INV_X32 U_g11954 ( .A(g11243), .ZN(g11954) );
INV_X32 U_g11958 ( .A(g11246), .ZN(g11958) );
INV_X32 U_g11959 ( .A(g11249), .ZN(g11959) );
INV_X32 U_g11960 ( .A(g11252), .ZN(g11960) );
INV_X32 U_g11961 ( .A(g11256), .ZN(g11961) );
INV_X32 U_g11963 ( .A(g11259), .ZN(g11963) );
INV_X32 U_g11968 ( .A(g11265), .ZN(g11968) );
INV_X32 U_g11969 ( .A(g11268), .ZN(g11969) );
INV_X32 U_g11970 ( .A(g11271), .ZN(g11970) );
INV_X32 U_g11971 ( .A(g11274), .ZN(g11971) );
INV_X32 U_g11972 ( .A(g11277), .ZN(g11972) );
INV_X32 U_g11973 ( .A(g11278), .ZN(g11973) );
INV_X32 U_I19160 ( .A(g10549), .ZN(I19160) );
INV_X32 U_g11976 ( .A(I19160), .ZN(g11976) );
INV_X32 U_g11982 ( .A(g11281), .ZN(g11982) );
INV_X32 U_g11983 ( .A(g11284), .ZN(g11983) );
INV_X32 U_g11984 ( .A(g11287), .ZN(g11984) );
INV_X32 U_g11985 ( .A(g11291), .ZN(g11985) );
INV_X32 U_g11986 ( .A(g11294), .ZN(g11986) );
INV_X32 U_g11989 ( .A(g11297), .ZN(g11989) );
INV_X32 U_I19174 ( .A(g9263), .ZN(I19174) );
INV_X32 U_g11990 ( .A(I19174), .ZN(g11990) );
INV_X32 U_g11994 ( .A(g11300), .ZN(g11994) );
INV_X32 U_g11995 ( .A(g11303), .ZN(g11995) );
INV_X32 U_g11996 ( .A(g11306), .ZN(g11996) );
INV_X32 U_g11997 ( .A(g11309), .ZN(g11997) );
INV_X32 U_g11998 ( .A(g11312), .ZN(g11998) );
INV_X32 U_g12001 ( .A(g11315), .ZN(g12001) );
INV_X32 U_g12002 ( .A(g11318), .ZN(g12002) );
INV_X32 U_g12003 ( .A(g11321), .ZN(g12003) );
INV_X32 U_g12004 ( .A(g11324), .ZN(g12004) );
INV_X32 U_g12007 ( .A(g11327), .ZN(g12007) );
INV_X32 U_I19195 ( .A(g8726), .ZN(I19195) );
INV_X32 U_g12009 ( .A(I19195), .ZN(g12009) );
INV_X32 U_g12013 ( .A(g10772), .ZN(g12013) );
INV_X32 U_g12017 ( .A(g10100), .ZN(g12017) );
INV_X32 U_g12020 ( .A(g11341), .ZN(g12020) );
INV_X32 U_g12021 ( .A(g11344), .ZN(g12021) );
INV_X32 U_g12022 ( .A(g11348), .ZN(g12022) );
INV_X32 U_g12023 ( .A(g11351), .ZN(g12023) );
INV_X32 U_g12024 ( .A(g11354), .ZN(g12024) );
INV_X32 U_g12025 ( .A(g11355), .ZN(g12025) );
INV_X32 U_I19208 ( .A(g10424), .ZN(I19208) );
INV_X32 U_g12027 ( .A(I19208), .ZN(g12027) );
INV_X32 U_I19211 ( .A(g10486), .ZN(I19211) );
INV_X32 U_g12030 ( .A(I19211), .ZN(g12030) );
INV_X32 U_g12037 ( .A(g11358), .ZN(g12037) );
INV_X32 U_g12038 ( .A(g11361), .ZN(g12038) );
INV_X32 U_g12039 ( .A(g11364), .ZN(g12039) );
INV_X32 U_g12040 ( .A(g11367), .ZN(g12040) );
INV_X32 U_g12041 ( .A(g11370), .ZN(g12041) );
INV_X32 U_g12042 ( .A(g11373), .ZN(g12042) );
INV_X32 U_I19226 ( .A(g10606), .ZN(I19226) );
INV_X32 U_g12045 ( .A(I19226), .ZN(g12045) );
INV_X32 U_g12051 ( .A(g11376), .ZN(g12051) );
INV_X32 U_g12052 ( .A(g11379), .ZN(g12052) );
INV_X32 U_g12053 ( .A(g11382), .ZN(g12053) );
INV_X32 U_g12054 ( .A(g11386), .ZN(g12054) );
INV_X32 U_g12055 ( .A(g11389), .ZN(g12055) );
INV_X32 U_g12058 ( .A(g11392), .ZN(g12058) );
INV_X32 U_I19240 ( .A(g9341), .ZN(I19240) );
INV_X32 U_g12059 ( .A(I19240), .ZN(g12059) );
INV_X32 U_g12063 ( .A(g11395), .ZN(g12063) );
INV_X32 U_g12064 ( .A(g11398), .ZN(g12064) );
INV_X32 U_g12065 ( .A(g11401), .ZN(g12065) );
INV_X32 U_g12066 ( .A(g11404), .ZN(g12066) );
INV_X32 U_g12067 ( .A(g11407), .ZN(g12067) );
INV_X32 U_g12071 ( .A(g10783), .ZN(g12071) );
INV_X32 U_g12075 ( .A(g11411), .ZN(g12075) );
INV_X32 U_g12076 ( .A(g11414), .ZN(g12076) );
INV_X32 U_g12077 ( .A(g11417), .ZN(g12077) );
INV_X32 U_g12078 ( .A(g11422), .ZN(g12078) );
INV_X32 U_g12084 ( .A(g11425), .ZN(g12084) );
INV_X32 U_g12085 ( .A(g11428), .ZN(g12085) );
INV_X32 U_g12086 ( .A(g11432), .ZN(g12086) );
INV_X32 U_g12087 ( .A(g11435), .ZN(g12087) );
INV_X32 U_g12088 ( .A(g11438), .ZN(g12088) );
INV_X32 U_g12089 ( .A(g11441), .ZN(g12089) );
INV_X32 U_I19271 ( .A(g10500), .ZN(I19271) );
INV_X32 U_g12091 ( .A(I19271), .ZN(g12091) );
INV_X32 U_I19274 ( .A(g10560), .ZN(I19274) );
INV_X32 U_g12094 ( .A(I19274), .ZN(g12094) );
INV_X32 U_g12101 ( .A(g11444), .ZN(g12101) );
INV_X32 U_g12102 ( .A(g11447), .ZN(g12102) );
INV_X32 U_g12103 ( .A(g11450), .ZN(g12103) );
INV_X32 U_g12104 ( .A(g11453), .ZN(g12104) );
INV_X32 U_g12105 ( .A(g11456), .ZN(g12105) );
INV_X32 U_g12106 ( .A(g11459), .ZN(g12106) );
INV_X32 U_I19289 ( .A(g10653), .ZN(I19289) );
INV_X32 U_g12109 ( .A(I19289), .ZN(g12109) );
INV_X32 U_g12115 ( .A(g11462), .ZN(g12115) );
INV_X32 U_g12116 ( .A(g11465), .ZN(g12116) );
INV_X32 U_g12117 ( .A(g11468), .ZN(g12117) );
INV_X32 U_g12118 ( .A(g11472), .ZN(g12118) );
INV_X32 U_g12119 ( .A(g11475), .ZN(g12119) );
INV_X32 U_g12122 ( .A(g11478), .ZN(g12122) );
INV_X32 U_I19303 ( .A(g9422), .ZN(I19303) );
INV_X32 U_g12123 ( .A(I19303), .ZN(g12123) );
INV_X32 U_I19307 ( .A(g8726), .ZN(I19307) );
INV_X32 U_g12125 ( .A(I19307), .ZN(g12125) );
INV_X32 U_g12130 ( .A(g10788), .ZN(g12130) );
INV_X32 U_g12134 ( .A(g8321), .ZN(g12134) );
INV_X32 U_g12135 ( .A(g8324), .ZN(g12135) );
INV_X32 U_I19315 ( .A(g10424), .ZN(I19315) );
INV_X32 U_g12136 ( .A(I19315), .ZN(g12136) );
INV_X32 U_I19318 ( .A(g10486), .ZN(I19318) );
INV_X32 U_g12139 ( .A(I19318), .ZN(g12139) );
INV_X32 U_I19321 ( .A(g10549), .ZN(I19321) );
INV_X32 U_g12142 ( .A(I19321), .ZN(g12142) );
INV_X32 U_g12147 ( .A(g8330), .ZN(g12147) );
INV_X32 U_g12148 ( .A(g8333), .ZN(g12148) );
INV_X32 U_g12149 ( .A(g8336), .ZN(g12149) );
INV_X32 U_g12150 ( .A(g8341), .ZN(g12150) );
INV_X32 U_g12156 ( .A(g8344), .ZN(g12156) );
INV_X32 U_g12157 ( .A(g8347), .ZN(g12157) );
INV_X32 U_g12158 ( .A(g8351), .ZN(g12158) );
INV_X32 U_g12159 ( .A(g8354), .ZN(g12159) );
INV_X32 U_g12160 ( .A(g8357), .ZN(g12160) );
INV_X32 U_g12161 ( .A(g8360), .ZN(g12161) );
INV_X32 U_I19342 ( .A(g10574), .ZN(I19342) );
INV_X32 U_g12163 ( .A(I19342), .ZN(g12163) );
INV_X32 U_I19345 ( .A(g10617), .ZN(I19345) );
INV_X32 U_g12166 ( .A(I19345), .ZN(g12166) );
INV_X32 U_g12173 ( .A(g8363), .ZN(g12173) );
INV_X32 U_g12174 ( .A(g8366), .ZN(g12174) );
INV_X32 U_g12175 ( .A(g8369), .ZN(g12175) );
INV_X32 U_g12176 ( .A(g8372), .ZN(g12176) );
INV_X32 U_g12177 ( .A(g8375), .ZN(g12177) );
INV_X32 U_g12178 ( .A(g8378), .ZN(g12178) );
INV_X32 U_I19360 ( .A(g10683), .ZN(I19360) );
INV_X32 U_g12181 ( .A(I19360), .ZN(g12181) );
INV_X32 U_g12187 ( .A(g8285), .ZN(g12187) );
INV_X32 U_g12191 ( .A(g8382), .ZN(g12191) );
INV_X32 U_g12196 ( .A(g8388), .ZN(g12196) );
INV_X32 U_g12197 ( .A(g8391), .ZN(g12197) );
INV_X32 U_I19374 ( .A(g10500), .ZN(I19374) );
INV_X32 U_g12198 ( .A(I19374), .ZN(g12198) );
INV_X32 U_I19377 ( .A(g10560), .ZN(I19377) );
INV_X32 U_g12201 ( .A(I19377), .ZN(g12201) );
INV_X32 U_I19380 ( .A(g10606), .ZN(I19380) );
INV_X32 U_g12204 ( .A(I19380), .ZN(g12204) );
INV_X32 U_g12209 ( .A(g8397), .ZN(g12209) );
INV_X32 U_g12210 ( .A(g8400), .ZN(g12210) );
INV_X32 U_g12211 ( .A(g8403), .ZN(g12211) );
INV_X32 U_g12212 ( .A(g8408), .ZN(g12212) );
INV_X32 U_g12218 ( .A(g8411), .ZN(g12218) );
INV_X32 U_g12219 ( .A(g8414), .ZN(g12219) );
INV_X32 U_g12220 ( .A(g8418), .ZN(g12220) );
INV_X32 U_g12221 ( .A(g8421), .ZN(g12221) );
INV_X32 U_g12222 ( .A(g8424), .ZN(g12222) );
INV_X32 U_g12223 ( .A(g8427), .ZN(g12223) );
INV_X32 U_I19401 ( .A(g10631), .ZN(I19401) );
INV_X32 U_g12225 ( .A(I19401), .ZN(g12225) );
INV_X32 U_I19404 ( .A(g10664), .ZN(I19404) );
INV_X32 U_g12228 ( .A(I19404), .ZN(g12228) );
INV_X32 U_g12235 ( .A(g8294), .ZN(g12235) );
INV_X32 U_I19412 ( .A(g10486), .ZN(I19412) );
INV_X32 U_g12239 ( .A(I19412), .ZN(g12239) );
INV_X32 U_I19415 ( .A(g10549), .ZN(I19415) );
INV_X32 U_g12242 ( .A(I19415), .ZN(g12242) );
INV_X32 U_g12246 ( .A(g8434), .ZN(g12246) );
INV_X32 U_g12251 ( .A(g8440), .ZN(g12251) );
INV_X32 U_g12252 ( .A(g8443), .ZN(g12252) );
INV_X32 U_I19426 ( .A(g10574), .ZN(I19426) );
INV_X32 U_g12253 ( .A(I19426), .ZN(g12253) );
INV_X32 U_I19429 ( .A(g10617), .ZN(I19429) );
INV_X32 U_g12256 ( .A(I19429), .ZN(g12256) );
INV_X32 U_I19432 ( .A(g10653), .ZN(I19432) );
INV_X32 U_g12259 ( .A(I19432), .ZN(g12259) );
INV_X32 U_g12264 ( .A(g8449), .ZN(g12264) );
INV_X32 U_g12265 ( .A(g8452), .ZN(g12265) );
INV_X32 U_g12266 ( .A(g8455), .ZN(g12266) );
INV_X32 U_g12267 ( .A(g8460), .ZN(g12267) );
INV_X32 U_g12275 ( .A(g8303), .ZN(g12275) );
INV_X32 U_I19449 ( .A(g10424), .ZN(I19449) );
INV_X32 U_g12279 ( .A(I19449), .ZN(g12279) );
INV_X32 U_I19452 ( .A(g10560), .ZN(I19452) );
INV_X32 U_g12282 ( .A(I19452), .ZN(g12282) );
INV_X32 U_I19455 ( .A(g10606), .ZN(I19455) );
INV_X32 U_g12285 ( .A(I19455), .ZN(g12285) );
INV_X32 U_g12289 ( .A(g8469), .ZN(g12289) );
INV_X32 U_g12294 ( .A(g8475), .ZN(g12294) );
INV_X32 U_g12295 ( .A(g8478), .ZN(g12295) );
INV_X32 U_I19466 ( .A(g10631), .ZN(I19466) );
INV_X32 U_g12296 ( .A(I19466), .ZN(g12296) );
INV_X32 U_I19469 ( .A(g10664), .ZN(I19469) );
INV_X32 U_g12299 ( .A(I19469), .ZN(g12299) );
INV_X32 U_I19472 ( .A(g10683), .ZN(I19472) );
INV_X32 U_g12302 ( .A(I19472), .ZN(g12302) );
INV_X32 U_g12308 ( .A(g8312), .ZN(g12308) );
INV_X32 U_I19479 ( .A(g10549), .ZN(I19479) );
INV_X32 U_g12312 ( .A(I19479), .ZN(g12312) );
INV_X32 U_I19482 ( .A(g10500), .ZN(I19482) );
INV_X32 U_g12315 ( .A(I19482), .ZN(g12315) );
INV_X32 U_I19485 ( .A(g10617), .ZN(I19485) );
INV_X32 U_g12318 ( .A(I19485), .ZN(g12318) );
INV_X32 U_I19488 ( .A(g10653), .ZN(I19488) );
INV_X32 U_g12321 ( .A(I19488), .ZN(g12321) );
INV_X32 U_g12325 ( .A(g8494), .ZN(g12325) );
INV_X32 U_g12332 ( .A(g10829), .ZN(g12332) );
INV_X32 U_I19500 ( .A(g10424), .ZN(I19500) );
INV_X32 U_g12333 ( .A(I19500), .ZN(g12333) );
INV_X32 U_I19503 ( .A(g10486), .ZN(I19503) );
INV_X32 U_g12336 ( .A(I19503), .ZN(g12336) );
INV_X32 U_I19507 ( .A(g10606), .ZN(I19507) );
INV_X32 U_g12340 ( .A(I19507), .ZN(g12340) );
INV_X32 U_I19510 ( .A(g10574), .ZN(I19510) );
INV_X32 U_g12343 ( .A(I19510), .ZN(g12343) );
INV_X32 U_I19513 ( .A(g10664), .ZN(I19513) );
INV_X32 U_g12346 ( .A(I19513), .ZN(g12346) );
INV_X32 U_I19516 ( .A(g10683), .ZN(I19516) );
INV_X32 U_g12349 ( .A(I19516), .ZN(g12349) );
INV_X32 U_g12354 ( .A(g8381), .ZN(g12354) );
INV_X32 U_g12362 ( .A(g10866), .ZN(g12362) );
INV_X32 U_I19523 ( .A(g10500), .ZN(I19523) );
INV_X32 U_g12363 ( .A(I19523), .ZN(g12363) );
INV_X32 U_I19526 ( .A(g10560), .ZN(I19526) );
INV_X32 U_g12366 ( .A(I19526), .ZN(g12366) );
INV_X32 U_I19530 ( .A(g10653), .ZN(I19530) );
INV_X32 U_g12370 ( .A(I19530), .ZN(g12370) );
INV_X32 U_I19533 ( .A(g10631), .ZN(I19533) );
INV_X32 U_g12373 ( .A(I19533), .ZN(g12373) );
INV_X32 U_g12378 ( .A(g10847), .ZN(g12378) );
INV_X32 U_I19539 ( .A(g10549), .ZN(I19539) );
INV_X32 U_g12379 ( .A(I19539), .ZN(g12379) );
INV_X32 U_I19542 ( .A(g10574), .ZN(I19542) );
INV_X32 U_g12382 ( .A(I19542), .ZN(g12382) );
INV_X32 U_I19545 ( .A(g10617), .ZN(I19545) );
INV_X32 U_g12385 ( .A(I19545), .ZN(g12385) );
INV_X32 U_I19549 ( .A(g10683), .ZN(I19549) );
INV_X32 U_g12389 ( .A(I19549), .ZN(g12389) );
INV_X32 U_I19552 ( .A(g8430), .ZN(I19552) );
INV_X32 U_g12392 ( .A(I19552), .ZN(g12392) );
INV_X32 U_g12408 ( .A(g11020), .ZN(g12408) );
INV_X32 U_I19557 ( .A(g10606), .ZN(I19557) );
INV_X32 U_g12409 ( .A(I19557), .ZN(g12409) );
INV_X32 U_I19560 ( .A(g10631), .ZN(I19560) );
INV_X32 U_g12412 ( .A(I19560), .ZN(g12412) );
INV_X32 U_I19563 ( .A(g10664), .ZN(I19563) );
INV_X32 U_g12415 ( .A(I19563), .ZN(g12415) );
INV_X32 U_g12420 ( .A(g10986), .ZN(g12420) );
INV_X32 U_I19569 ( .A(g10653), .ZN(I19569) );
INV_X32 U_g12421 ( .A(I19569), .ZN(g12421) );
INV_X32 U_g12424 ( .A(g10962), .ZN(g12424) );
INV_X32 U_I19573 ( .A(g8835), .ZN(I19573) );
INV_X32 U_g12425 ( .A(I19573), .ZN(g12425) );
INV_X32 U_I19576 ( .A(g10683), .ZN(I19576) );
INV_X32 U_g12426 ( .A(I19576), .ZN(g12426) );
INV_X32 U_g12430 ( .A(g10905), .ZN(g12430) );
INV_X32 U_I19582 ( .A(g8862), .ZN(I19582) );
INV_X32 U_g12432 ( .A(I19582), .ZN(g12432) );
INV_X32 U_g12434 ( .A(g10929), .ZN(g12434) );
INV_X32 U_I19587 ( .A(g9173), .ZN(I19587) );
INV_X32 U_g12435 ( .A(I19587), .ZN(g12435) );
INV_X32 U_I19591 ( .A(g8900), .ZN(I19591) );
INV_X32 U_g12437 ( .A(I19591), .ZN(g12437) );
INV_X32 U_g12438 ( .A(g10846), .ZN(g12438) );
INV_X32 U_I19595 ( .A(g10810), .ZN(I19595) );
INV_X32 U_g12439 ( .A(I19595), .ZN(g12439) );
INV_X32 U_I19598 ( .A(g9215), .ZN(I19598) );
INV_X32 U_g12440 ( .A(I19598), .ZN(g12440) );
INV_X32 U_I19602 ( .A(g8940), .ZN(I19602) );
INV_X32 U_g12442 ( .A(I19602), .ZN(g12442) );
INV_X32 U_I19605 ( .A(g10797), .ZN(I19605) );
INV_X32 U_g12443 ( .A(I19605), .ZN(g12443) );
INV_X32 U_I19608 ( .A(g10831), .ZN(I19608) );
INV_X32 U_g12444 ( .A(I19608), .ZN(g12444) );
INV_X32 U_I19611 ( .A(g9276), .ZN(I19611) );
INV_X32 U_g12445 ( .A(I19611), .ZN(g12445) );
INV_X32 U_I19615 ( .A(g10789), .ZN(I19615) );
INV_X32 U_g12447 ( .A(I19615), .ZN(g12447) );
INV_X32 U_I19618 ( .A(g10814), .ZN(I19618) );
INV_X32 U_g12448 ( .A(I19618), .ZN(g12448) );
INV_X32 U_I19621 ( .A(g10851), .ZN(I19621) );
INV_X32 U_g12449 ( .A(I19621), .ZN(g12449) );
INV_X32 U_I19624 ( .A(g9354), .ZN(I19624) );
INV_X32 U_g12450 ( .A(I19624), .ZN(g12450) );
INV_X32 U_I19628 ( .A(g10784), .ZN(I19628) );
INV_X32 U_g12452 ( .A(I19628), .ZN(g12452) );
INV_X32 U_I19631 ( .A(g10801), .ZN(I19631) );
INV_X32 U_g12453 ( .A(I19631), .ZN(g12453) );
INV_X32 U_I19634 ( .A(g10835), .ZN(I19634) );
INV_X32 U_g12454 ( .A(I19634), .ZN(g12454) );
INV_X32 U_I19637 ( .A(g10872), .ZN(I19637) );
INV_X32 U_g12455 ( .A(I19637), .ZN(g12455) );
INV_X32 U_g12456 ( .A(g8602), .ZN(g12456) );
INV_X32 U_I19642 ( .A(g10793), .ZN(I19642) );
INV_X32 U_g12460 ( .A(I19642), .ZN(g12460) );
INV_X32 U_I19645 ( .A(g10818), .ZN(I19645) );
INV_X32 U_g12461 ( .A(I19645), .ZN(g12461) );
INV_X32 U_I19648 ( .A(g10855), .ZN(I19648) );
INV_X32 U_g12462 ( .A(I19648), .ZN(g12462) );
INV_X32 U_g12463 ( .A(g10730), .ZN(g12463) );
INV_X32 U_g12466 ( .A(g8614), .ZN(g12466) );
INV_X32 U_I19654 ( .A(g10805), .ZN(I19654) );
INV_X32 U_g12470 ( .A(I19654), .ZN(g12470) );
INV_X32 U_I19657 ( .A(g10839), .ZN(I19657) );
INV_X32 U_g12471 ( .A(I19657), .ZN(g12471) );
INV_X32 U_g12472 ( .A(g8617), .ZN(g12472) );
INV_X32 U_g12473 ( .A(g8580), .ZN(g12473) );
INV_X32 U_g12476 ( .A(g8622), .ZN(g12476) );
INV_X32 U_g12478 ( .A(g10749), .ZN(g12478) );
INV_X32 U_g12481 ( .A(g8627), .ZN(g12481) );
INV_X32 U_I19667 ( .A(g10822), .ZN(I19667) );
INV_X32 U_g12485 ( .A(I19667), .ZN(g12485) );
INV_X32 U_g12490 ( .A(g8587), .ZN(g12490) );
INV_X32 U_g12493 ( .A(g8632), .ZN(g12493) );
INV_X32 U_g12495 ( .A(g10767), .ZN(g12495) );
INV_X32 U_g12498 ( .A(g8637), .ZN(g12498) );
INV_X32 U_g12502 ( .A(g8640), .ZN(g12502) );
INV_X32 U_g12504 ( .A(g8643), .ZN(g12504) );
INV_X32 U_g12505 ( .A(g8646), .ZN(g12505) );
INV_X32 U_g12510 ( .A(g8594), .ZN(g12510) );
INV_X32 U_g12513 ( .A(g8651), .ZN(g12513) );
INV_X32 U_g12515 ( .A(g10773), .ZN(g12515) );
INV_X32 U_g12518 ( .A(g8655), .ZN(g12518) );
INV_X32 U_I19689 ( .A(g10016), .ZN(I19689) );
INV_X32 U_g12519 ( .A(I19689), .ZN(g12519) );
INV_X32 U_g12521 ( .A(g8659), .ZN(g12521) );
INV_X32 U_g12522 ( .A(g8662), .ZN(g12522) );
INV_X32 U_g12527 ( .A(g8605), .ZN(g12527) );
INV_X32 U_g12530 ( .A(g8667), .ZN(g12530) );
INV_X32 U_g12532 ( .A(g8670), .ZN(g12532) );
INV_X32 U_g12533 ( .A(g8673), .ZN(g12533) );
INV_X32 U_I19702 ( .A(g10125), .ZN(I19702) );
INV_X32 U_g12534 ( .A(I19702), .ZN(g12534) );
INV_X32 U_g12536 ( .A(g8678), .ZN(g12536) );
INV_X32 U_g12537 ( .A(g8681), .ZN(g12537) );
INV_X32 U_g12542 ( .A(g8684), .ZN(g12542) );
INV_X32 U_I19711 ( .A(g10230), .ZN(I19711) );
INV_X32 U_g12543 ( .A(I19711), .ZN(g12543) );
INV_X32 U_g12545 ( .A(g8690), .ZN(g12545) );
INV_X32 U_g12546 ( .A(g8693), .ZN(g12546) );
INV_X32 U_g12547 ( .A(g8696), .ZN(g12547) );
INV_X32 U_I19718 ( .A(g8726), .ZN(I19718) );
INV_X32 U_g12548 ( .A(I19718), .ZN(g12548) );
INV_X32 U_g12551 ( .A(g8700), .ZN(g12551) );
INV_X32 U_I19722 ( .A(g10332), .ZN(I19722) );
INV_X32 U_g12552 ( .A(I19722), .ZN(g12552) );
INV_X32 U_g12553 ( .A(g8708), .ZN(g12553) );
INV_X32 U_g12554 ( .A(g8711), .ZN(g12554) );
INV_X32 U_I19727 ( .A(g8726), .ZN(I19727) );
INV_X32 U_g12555 ( .A(I19727), .ZN(g12555) );
INV_X32 U_g12558 ( .A(g8714), .ZN(g12558) );
INV_X32 U_g12559 ( .A(g8719), .ZN(g12559) );
INV_X32 U_g12560 ( .A(g8745), .ZN(g12560) );
INV_X32 U_I19733 ( .A(g8726), .ZN(I19733) );
INV_X32 U_g12561 ( .A(I19733), .ZN(g12561) );
INV_X32 U_I19736 ( .A(g9184), .ZN(I19736) );
INV_X32 U_g12564 ( .A(I19736), .ZN(g12564) );
INV_X32 U_I19739 ( .A(g10694), .ZN(I19739) );
INV_X32 U_g12565 ( .A(I19739), .ZN(g12565) );
INV_X32 U_g12596 ( .A(g8748), .ZN(g12596) );
INV_X32 U_g12597 ( .A(g8752), .ZN(g12597) );
INV_X32 U_g12598 ( .A(g8757), .ZN(g12598) );
INV_X32 U_g12599 ( .A(g8763), .ZN(g12599) );
INV_X32 U_g12600 ( .A(g8766), .ZN(g12600) );
INV_X32 U_I19747 ( .A(g8726), .ZN(I19747) );
INV_X32 U_g12601 ( .A(I19747), .ZN(g12601) );
INV_X32 U_I19750 ( .A(g8726), .ZN(I19750) );
INV_X32 U_g12604 ( .A(I19750), .ZN(g12604) );
INV_X32 U_I19753 ( .A(g9229), .ZN(I19753) );
INV_X32 U_g12607 ( .A(I19753), .ZN(g12607) );
INV_X32 U_I19756 ( .A(g10424), .ZN(I19756) );
INV_X32 U_g12608 ( .A(I19756), .ZN(g12608) );
INV_X32 U_I19759 ( .A(g10714), .ZN(I19759) );
INV_X32 U_g12611 ( .A(I19759), .ZN(g12611) );
INV_X32 U_g12642 ( .A(g8771), .ZN(g12642) );
INV_X32 U_g12643 ( .A(g8775), .ZN(g12643) );
INV_X32 U_g12644 ( .A(g8780), .ZN(g12644) );
INV_X32 U_g12645 ( .A(g8785), .ZN(g12645) );
INV_X32 U_g12646 ( .A(g8788), .ZN(g12646) );
INV_X32 U_I19767 ( .A(g8726), .ZN(I19767) );
INV_X32 U_g12647 ( .A(I19767), .ZN(g12647) );
INV_X32 U_I19771 ( .A(g10038), .ZN(I19771) );
INV_X32 U_g12651 ( .A(I19771), .ZN(g12651) );
INV_X32 U_I19774 ( .A(g10500), .ZN(I19774) );
INV_X32 U_g12654 ( .A(I19774), .ZN(g12654) );
INV_X32 U_I19777 ( .A(g10735), .ZN(I19777) );
INV_X32 U_g12657 ( .A(I19777), .ZN(g12657) );
INV_X32 U_g12688 ( .A(g8794), .ZN(g12688) );
INV_X32 U_g12689 ( .A(g8798), .ZN(g12689) );
INV_X32 U_g12690 ( .A(g8802), .ZN(g12690) );
INV_X32 U_g12691 ( .A(g8805), .ZN(g12691) );
INV_X32 U_I19784 ( .A(g8726), .ZN(I19784) );
INV_X32 U_g12692 ( .A(I19784), .ZN(g12692) );
INV_X32 U_I19787 ( .A(g8726), .ZN(I19787) );
INV_X32 U_g12695 ( .A(I19787), .ZN(g12695) );
INV_X32 U_I19791 ( .A(g10486), .ZN(I19791) );
INV_X32 U_g12699 ( .A(I19791), .ZN(g12699) );
INV_X32 U_I19794 ( .A(g10676), .ZN(I19794) );
INV_X32 U_g12702 ( .A(I19794), .ZN(g12702) );
INV_X32 U_I19797 ( .A(g10147), .ZN(I19797) );
INV_X32 U_g12705 ( .A(I19797), .ZN(g12705) );
INV_X32 U_I19800 ( .A(g10574), .ZN(I19800) );
INV_X32 U_g12708 ( .A(I19800), .ZN(g12708) );
INV_X32 U_I19803 ( .A(g10754), .ZN(I19803) );
INV_X32 U_g12711 ( .A(I19803), .ZN(g12711) );
INV_X32 U_g12742 ( .A(g8813), .ZN(g12742) );
INV_X32 U_g12743 ( .A(g8817), .ZN(g12743) );
INV_X32 U_I19808 ( .A(g8726), .ZN(I19808) );
INV_X32 U_g12744 ( .A(I19808), .ZN(g12744) );
INV_X32 U_g12748 ( .A(g8823), .ZN(g12748) );
INV_X32 U_I19813 ( .A(g10649), .ZN(I19813) );
INV_X32 U_g12749 ( .A(I19813), .ZN(g12749) );
INV_X32 U_I19816 ( .A(g10703), .ZN(I19816) );
INV_X32 U_g12752 ( .A(I19816), .ZN(g12752) );
INV_X32 U_I19820 ( .A(g10560), .ZN(I19820) );
INV_X32 U_g12756 ( .A(I19820), .ZN(g12756) );
INV_X32 U_I19823 ( .A(g10705), .ZN(I19823) );
INV_X32 U_g12759 ( .A(I19823), .ZN(g12759) );
INV_X32 U_I19826 ( .A(g10252), .ZN(I19826) );
INV_X32 U_g12762 ( .A(I19826), .ZN(g12762) );
INV_X32 U_I19829 ( .A(g10631), .ZN(I19829) );
INV_X32 U_g12765 ( .A(I19829), .ZN(g12765) );
INV_X32 U_g12768 ( .A(g8829), .ZN(g12768) );
INV_X32 U_I19833 ( .A(g8726), .ZN(I19833) );
INV_X32 U_g12769 ( .A(I19833), .ZN(g12769) );
INV_X32 U_I19836 ( .A(g8726), .ZN(I19836) );
INV_X32 U_g12772 ( .A(I19836), .ZN(g12772) );
INV_X32 U_g12775 ( .A(g8832), .ZN(g12775) );
INV_X32 U_g12776 ( .A(g10766), .ZN(g12776) );
INV_X32 U_g12782 ( .A(g8836), .ZN(g12782) );
INV_X32 U_I19844 ( .A(g8533), .ZN(I19844) );
INV_X32 U_g12783 ( .A(I19844), .ZN(g12783) );
INV_X32 U_I19847 ( .A(g10677), .ZN(I19847) );
INV_X32 U_g12786 ( .A(I19847), .ZN(g12786) );
INV_X32 U_g12790 ( .A(g8847), .ZN(g12790) );
INV_X32 U_I19852 ( .A(g10679), .ZN(I19852) );
INV_X32 U_g12791 ( .A(I19852), .ZN(g12791) );
INV_X32 U_I19855 ( .A(g10723), .ZN(I19855) );
INV_X32 U_g12794 ( .A(I19855), .ZN(g12794) );
INV_X32 U_I19859 ( .A(g10617), .ZN(I19859) );
INV_X32 U_g12798 ( .A(I19859), .ZN(g12798) );
INV_X32 U_I19862 ( .A(g10725), .ZN(I19862) );
INV_X32 U_g12801 ( .A(I19862), .ZN(g12801) );
INV_X32 U_I19865 ( .A(g10354), .ZN(I19865) );
INV_X32 U_g12804 ( .A(I19865), .ZN(g12804) );
INV_X32 U_g12807 ( .A(g8853), .ZN(g12807) );
INV_X32 U_I19869 ( .A(g8726), .ZN(I19869) );
INV_X32 U_g12808 ( .A(I19869), .ZN(g12808) );
INV_X32 U_I19872 ( .A(g8317), .ZN(I19872) );
INV_X32 U_g12811 ( .A(I19872), .ZN(g12811) );
INV_X32 U_g12815 ( .A(g8856), .ZN(g12815) );
INV_X32 U_I19877 ( .A(g8547), .ZN(I19877) );
INV_X32 U_g12816 ( .A(I19877), .ZN(g12816) );
INV_X32 U_g12821 ( .A(g8863), .ZN(g12821) );
INV_X32 U_I19883 ( .A(g8550), .ZN(I19883) );
INV_X32 U_g12822 ( .A(I19883), .ZN(g12822) );
INV_X32 U_I19886 ( .A(g10706), .ZN(I19886) );
INV_X32 U_g12825 ( .A(I19886), .ZN(g12825) );
INV_X32 U_g12829 ( .A(g8874), .ZN(g12829) );
INV_X32 U_I19891 ( .A(g10708), .ZN(I19891) );
INV_X32 U_g12830 ( .A(I19891), .ZN(g12830) );
INV_X32 U_I19894 ( .A(g10744), .ZN(I19894) );
INV_X32 U_g12833 ( .A(I19894), .ZN(g12833) );
INV_X32 U_I19898 ( .A(g10664), .ZN(I19898) );
INV_X32 U_g12837 ( .A(I19898), .ZN(g12837) );
INV_X32 U_I19901 ( .A(g10746), .ZN(I19901) );
INV_X32 U_g12840 ( .A(I19901), .ZN(g12840) );
INV_X32 U_g12843 ( .A(g8879), .ZN(g12843) );
INV_X32 U_I19905 ( .A(g8726), .ZN(I19905) );
INV_X32 U_g12844 ( .A(I19905), .ZN(g12844) );
INV_X32 U_g12847 ( .A(g8882), .ZN(g12847) );
INV_X32 U_g12848 ( .A(g11059), .ZN(g12848) );
INV_X32 U_g12850 ( .A(g8885), .ZN(g12850) );
INV_X32 U_g12851 ( .A(g8888), .ZN(g12851) );
INV_X32 U_g12853 ( .A(g8894), .ZN(g12853) );
INV_X32 U_I19915 ( .A(g8560), .ZN(I19915) );
INV_X32 U_g12854 ( .A(I19915), .ZN(g12854) );
INV_X32 U_g12859 ( .A(g8901), .ZN(g12859) );
INV_X32 U_I19921 ( .A(g8563), .ZN(I19921) );
INV_X32 U_g12860 ( .A(I19921), .ZN(g12860) );
INV_X32 U_I19924 ( .A(g10726), .ZN(I19924) );
INV_X32 U_g12863 ( .A(I19924), .ZN(g12863) );
INV_X32 U_g12867 ( .A(g8912), .ZN(g12867) );
INV_X32 U_I19929 ( .A(g10728), .ZN(I19929) );
INV_X32 U_g12868 ( .A(I19929), .ZN(g12868) );
INV_X32 U_I19932 ( .A(g10763), .ZN(I19932) );
INV_X32 U_g12871 ( .A(I19932), .ZN(g12871) );
INV_X32 U_g12874 ( .A(g8915), .ZN(g12874) );
INV_X32 U_g12875 ( .A(g10779), .ZN(g12875) );
INV_X32 U_g12881 ( .A(g8918), .ZN(g12881) );
INV_X32 U_g12882 ( .A(g8921), .ZN(g12882) );
INV_X32 U_g12891 ( .A(g8925), .ZN(g12891) );
INV_X32 U_g12892 ( .A(g8928), .ZN(g12892) );
INV_X32 U_g12894 ( .A(g8934), .ZN(g12894) );
INV_X32 U_I19952 ( .A(g8571), .ZN(I19952) );
INV_X32 U_g12895 ( .A(I19952), .ZN(g12895) );
INV_X32 U_g12900 ( .A(g8941), .ZN(g12900) );
INV_X32 U_I19958 ( .A(g8574), .ZN(I19958) );
INV_X32 U_g12901 ( .A(I19958), .ZN(g12901) );
INV_X32 U_I19961 ( .A(g10747), .ZN(I19961) );
INV_X32 U_g12904 ( .A(I19961), .ZN(g12904) );
INV_X32 U_g12907 ( .A(g8949), .ZN(g12907) );
INV_X32 U_g12909 ( .A(g10904), .ZN(g12909) );
INV_X32 U_g12914 ( .A(g8952), .ZN(g12914) );
INV_X32 U_g12915 ( .A(g8955), .ZN(g12915) );
INV_X32 U_g12921 ( .A(g8958), .ZN(g12921) );
INV_X32 U_g12922 ( .A(g8961), .ZN(g12922) );
INV_X32 U_g12931 ( .A(g8965), .ZN(g12931) );
INV_X32 U_g12932 ( .A(g8968), .ZN(g12932) );
INV_X32 U_g12934 ( .A(g8974), .ZN(g12934) );
INV_X32 U_I19986 ( .A(g8577), .ZN(I19986) );
INV_X32 U_g12935 ( .A(I19986), .ZN(g12935) );
INV_X32 U_g12940 ( .A(g8980), .ZN(g12940) );
INV_X32 U_g12943 ( .A(g8984), .ZN(g12943) );
INV_X32 U_g12944 ( .A(g8987), .ZN(g12944) );
INV_X32 U_g12950 ( .A(g8990), .ZN(g12950) );
INV_X32 U_g12951 ( .A(g8993), .ZN(g12951) );
INV_X32 U_g12960 ( .A(g8997), .ZN(g12960) );
INV_X32 U_g12961 ( .A(g9000), .ZN(g12961) );
INV_X32 U_I20009 ( .A(g8313), .ZN(I20009) );
INV_X32 U_g12962 ( .A(I20009), .ZN(g12962) );
INV_X32 U_g12965 ( .A(g9006), .ZN(g12965) );
INV_X32 U_g12969 ( .A(g9010), .ZN(g12969) );
INV_X32 U_g12972 ( .A(g9013), .ZN(g12972) );
INV_X32 U_g12973 ( .A(g9016), .ZN(g12973) );
INV_X32 U_g12979 ( .A(g9019), .ZN(g12979) );
INV_X32 U_g12980 ( .A(g9022), .ZN(g12980) );
INV_X32 U_g12993 ( .A(g9035), .ZN(g12993) );
INV_X32 U_g12996 ( .A(g9038), .ZN(g12996) );
INV_X32 U_g12997 ( .A(g9041), .ZN(g12997) );
INV_X32 U_g12998 ( .A(g9044), .ZN(g12998) );
INV_X32 U_g13003 ( .A(g9058), .ZN(g13003) );
INV_X32 U_I20062 ( .A(g10480), .ZN(I20062) );
INV_X32 U_g13011 ( .A(I20062), .ZN(g13011) );
INV_X32 U_g13025 ( .A(g10810), .ZN(g13025) );
INV_X32 U_g13033 ( .A(g10797), .ZN(g13033) );
INV_X32 U_g13036 ( .A(g10831), .ZN(g13036) );
INV_X32 U_g13043 ( .A(g10789), .ZN(g13043) );
INV_X32 U_g13046 ( .A(g10814), .ZN(g13046) );
INV_X32 U_g13049 ( .A(g10851), .ZN(g13049) );
INV_X32 U_g13057 ( .A(g10784), .ZN(g13057) );
INV_X32 U_g13060 ( .A(g10801), .ZN(g13060) );
INV_X32 U_g13063 ( .A(g10835), .ZN(g13063) );
INV_X32 U_g13066 ( .A(g10872), .ZN(g13066) );
INV_X32 U_I20117 ( .A(g10876), .ZN(I20117) );
INV_X32 U_g13070 ( .A(I20117), .ZN(g13070) );
INV_X32 U_g13073 ( .A(g10793), .ZN(g13073) );
INV_X32 U_g13076 ( .A(g10818), .ZN(g13076) );
INV_X32 U_g13079 ( .A(g10855), .ZN(g13079) );
INV_X32 U_g13092 ( .A(g10805), .ZN(g13092) );
INV_X32 U_g13095 ( .A(g10839), .ZN(g13095) );
INV_X32 U_g13101 ( .A(g9128), .ZN(g13101) );
INV_X32 U_g13107 ( .A(g10822), .ZN(g13107) );
INV_X32 U_g13117 ( .A(g9134), .ZN(g13117) );
INV_X32 U_g13130 ( .A(g9140), .ZN(g13130) );
INV_X32 U_g13141 ( .A(g9146), .ZN(g13141) );
INV_X32 U_g13148 ( .A(g9170), .ZN(g13148) );
INV_X32 U_g13151 ( .A(g9184), .ZN(g13151) );
INV_X32 U_g13152 ( .A(g9196), .ZN(g13152) );
INV_X32 U_g13153 ( .A(g9199), .ZN(g13153) );
INV_X32 U_g13154 ( .A(g9212), .ZN(g13154) );
INV_X32 U_g13157 ( .A(g9229), .ZN(g13157) );
INV_X32 U_g13158 ( .A(g9242), .ZN(g13158) );
INV_X32 U_g13159 ( .A(g9245), .ZN(g13159) );
INV_X32 U_g13161 ( .A(g9257), .ZN(g13161) );
INV_X32 U_g13162 ( .A(g9260), .ZN(g13162) );
INV_X32 U_g13163 ( .A(g9273), .ZN(g13163) );
INV_X32 U_g13166 ( .A(g9290), .ZN(g13166) );
INV_X32 U_g13167 ( .A(g9303), .ZN(g13167) );
INV_X32 U_g13168 ( .A(g9306), .ZN(g13168) );
INV_X32 U_g13169 ( .A(g9320), .ZN(g13169) );
INV_X32 U_g13170 ( .A(g9323), .ZN(g13170) );
INV_X32 U_g13172 ( .A(g9335), .ZN(g13172) );
INV_X32 U_g13173 ( .A(g9338), .ZN(g13173) );
INV_X32 U_g13174 ( .A(g9351), .ZN(g13174) );
INV_X32 U_g13176 ( .A(g9368), .ZN(g13176) );
INV_X32 U_g13177 ( .A(g9371), .ZN(g13177) );
INV_X32 U_g13178 ( .A(g9384), .ZN(g13178) );
INV_X32 U_g13179 ( .A(g9387), .ZN(g13179) );
INV_X32 U_g13180 ( .A(g9401), .ZN(g13180) );
INV_X32 U_g13181 ( .A(g9404), .ZN(g13181) );
INV_X32 U_g13183 ( .A(g9416), .ZN(g13183) );
INV_X32 U_g13184 ( .A(g9419), .ZN(g13184) );
INV_X32 U_g13185 ( .A(g9443), .ZN(g13185) );
INV_X32 U_g13186 ( .A(g9446), .ZN(g13186) );
INV_X32 U_g13187 ( .A(g9450), .ZN(g13187) );
INV_X32 U_g13188 ( .A(g9465), .ZN(g13188) );
INV_X32 U_g13189 ( .A(g9468), .ZN(g13189) );
INV_X32 U_g13190 ( .A(g9481), .ZN(g13190) );
INV_X32 U_g13191 ( .A(g9484), .ZN(g13191) );
INV_X32 U_g13192 ( .A(g9498), .ZN(g13192) );
INV_X32 U_g13193 ( .A(g9501), .ZN(g13193) );
INV_X32 U_g13195 ( .A(g9524), .ZN(g13195) );
INV_X32 U_g13196 ( .A(g9528), .ZN(g13196) );
INV_X32 U_g13197 ( .A(g9531), .ZN(g13197) );
INV_X32 U_g13198 ( .A(g9585), .ZN(g13198) );
INV_X32 U_g13199 ( .A(g9588), .ZN(g13199) );
INV_X32 U_g13200 ( .A(g9592), .ZN(g13200) );
INV_X32 U_g13201 ( .A(g9607), .ZN(g13201) );
INV_X32 U_g13202 ( .A(g9610), .ZN(g13202) );
INV_X32 U_g13203 ( .A(g9623), .ZN(g13203) );
INV_X32 U_g13204 ( .A(g9626), .ZN(g13204) );
INV_X32 U_g13205 ( .A(g9641), .ZN(g13205) );
INV_X32 U_g13206 ( .A(g9644), .ZN(g13206) );
INV_X32 U_g13207 ( .A(g9666), .ZN(g13207) );
INV_X32 U_g13208 ( .A(g9670), .ZN(g13208) );
INV_X32 U_g13209 ( .A(g9673), .ZN(g13209) );
INV_X32 U_g13210 ( .A(g9727), .ZN(g13210) );
INV_X32 U_g13211 ( .A(g9730), .ZN(g13211) );
INV_X32 U_g13212 ( .A(g9734), .ZN(g13212) );
INV_X32 U_g13213 ( .A(g9749), .ZN(g13213) );
INV_X32 U_g13214 ( .A(g9752), .ZN(g13214) );
INV_X32 U_I20264 ( .A(g9027), .ZN(I20264) );
INV_X32 U_g13215 ( .A(I20264), .ZN(g13215) );
INV_X32 U_g13218 ( .A(g9767), .ZN(g13218) );
INV_X32 U_g13219 ( .A(g9770), .ZN(g13219) );
INV_X32 U_g13220 ( .A(g9787), .ZN(g13220) );
INV_X32 U_g13221 ( .A(g9790), .ZN(g13221) );
INV_X32 U_g13222 ( .A(g9812), .ZN(g13222) );
INV_X32 U_g13223 ( .A(g9816), .ZN(g13223) );
INV_X32 U_g13224 ( .A(g9819), .ZN(g13224) );
INV_X32 U_g13225 ( .A(g9873), .ZN(g13225) );
INV_X32 U_g13226 ( .A(g9876), .ZN(g13226) );
INV_X32 U_g13227 ( .A(g9880), .ZN(g13227) );
INV_X32 U_I20278 ( .A(g9027), .ZN(I20278) );
INV_X32 U_g13229 ( .A(I20278), .ZN(g13229) );
INV_X32 U_g13232 ( .A(g9895), .ZN(g13232) );
INV_X32 U_g13233 ( .A(g9898), .ZN(g13233) );
INV_X32 U_I20283 ( .A(g9050), .ZN(I20283) );
INV_X32 U_g13234 ( .A(I20283), .ZN(g13234) );
INV_X32 U_g13237 ( .A(g9913), .ZN(g13237) );
INV_X32 U_g13238 ( .A(g9916), .ZN(g13238) );
INV_X32 U_g13239 ( .A(g9933), .ZN(g13239) );
INV_X32 U_g13240 ( .A(g9936), .ZN(g13240) );
INV_X32 U_g13241 ( .A(g9958), .ZN(g13241) );
INV_X32 U_g13242 ( .A(g9962), .ZN(g13242) );
INV_X32 U_g13243 ( .A(g9965), .ZN(g13243) );
INV_X32 U_g13244 ( .A(g10004), .ZN(g13244) );
INV_X32 U_I20295 ( .A(g10015), .ZN(I20295) );
INV_X32 U_g13246 ( .A(I20295), .ZN(g13246) );
INV_X32 U_I20299 ( .A(g10800), .ZN(I20299) );
INV_X32 U_g13248 ( .A(I20299), .ZN(g13248) );
INV_X32 U_g13249 ( .A(g10018), .ZN(g13249) );
INV_X32 U_g13250 ( .A(g10021), .ZN(g13250) );
INV_X32 U_I20305 ( .A(g9050), .ZN(I20305) );
INV_X32 U_g13252 ( .A(I20305), .ZN(g13252) );
INV_X32 U_g13255 ( .A(g10049), .ZN(g13255) );
INV_X32 U_g13256 ( .A(g10052), .ZN(g13256) );
INV_X32 U_I20310 ( .A(g9067), .ZN(I20310) );
INV_X32 U_g13257 ( .A(I20310), .ZN(g13257) );
INV_X32 U_g13260 ( .A(g10067), .ZN(g13260) );
INV_X32 U_g13261 ( .A(g10070), .ZN(g13261) );
INV_X32 U_g13262 ( .A(g10087), .ZN(g13262) );
INV_X32 U_g13263 ( .A(g10090), .ZN(g13263) );
INV_X32 U_g13264 ( .A(g10096), .ZN(g13264) );
INV_X32 U_g13265 ( .A(g8568), .ZN(g13265) );
INV_X32 U_I20320 ( .A(g10792), .ZN(I20320) );
INV_X32 U_g13267 ( .A(I20320), .ZN(g13267) );
INV_X32 U_g13268 ( .A(g10109), .ZN(g13268) );
INV_X32 U_I20324 ( .A(g10124), .ZN(I20324) );
INV_X32 U_g13269 ( .A(I20324), .ZN(g13269) );
INV_X32 U_I20328 ( .A(g10817), .ZN(I20328) );
INV_X32 U_g13271 ( .A(I20328), .ZN(g13271) );
INV_X32 U_g13272 ( .A(g10127), .ZN(g13272) );
INV_X32 U_g13273 ( .A(g10130), .ZN(g13273) );
INV_X32 U_I20334 ( .A(g9067), .ZN(I20334) );
INV_X32 U_g13275 ( .A(I20334), .ZN(g13275) );
INV_X32 U_g13278 ( .A(g10158), .ZN(g13278) );
INV_X32 U_g13279 ( .A(g10161), .ZN(g13279) );
INV_X32 U_I20339 ( .A(g9084), .ZN(I20339) );
INV_X32 U_g13280 ( .A(I20339), .ZN(g13280) );
INV_X32 U_g13283 ( .A(g10176), .ZN(g13283) );
INV_X32 U_g13284 ( .A(g10179), .ZN(g13284) );
INV_X32 U_g13285 ( .A(g10189), .ZN(g13285) );
INV_X32 U_I20347 ( .A(g10787), .ZN(I20347) );
INV_X32 U_g13290 ( .A(I20347), .ZN(g13290) );
INV_X32 U_I20351 ( .A(g10804), .ZN(I20351) );
INV_X32 U_g13292 ( .A(I20351), .ZN(g13292) );
INV_X32 U_g13293 ( .A(g10214), .ZN(g13293) );
INV_X32 U_I20355 ( .A(g10229), .ZN(I20355) );
INV_X32 U_g13294 ( .A(I20355), .ZN(g13294) );
INV_X32 U_I20359 ( .A(g10838), .ZN(I20359) );
INV_X32 U_g13296 ( .A(I20359), .ZN(g13296) );
INV_X32 U_g13297 ( .A(g10232), .ZN(g13297) );
INV_X32 U_g13298 ( .A(g10235), .ZN(g13298) );
INV_X32 U_I20365 ( .A(g9084), .ZN(I20365) );
INV_X32 U_g13300 ( .A(I20365), .ZN(g13300) );
INV_X32 U_g13303 ( .A(g10263), .ZN(g13303) );
INV_X32 U_g13304 ( .A(g10266), .ZN(g13304) );
INV_X32 U_g13308 ( .A(g10273), .ZN(g13308) );
INV_X32 U_g13309 ( .A(g10276), .ZN(g13309) );
INV_X32 U_I20376 ( .A(g8569), .ZN(I20376) );
INV_X32 U_g13317 ( .A(I20376), .ZN(g13317) );
INV_X32 U_I20379 ( .A(g11213), .ZN(I20379) );
INV_X32 U_g13318 ( .A(I20379), .ZN(g13318) );
INV_X32 U_I20382 ( .A(g10907), .ZN(I20382) );
INV_X32 U_g13319 ( .A(I20382), .ZN(g13319) );
INV_X32 U_I20386 ( .A(g10796), .ZN(I20386) );
INV_X32 U_g13321 ( .A(I20386), .ZN(g13321) );
INV_X32 U_I20390 ( .A(g10821), .ZN(I20390) );
INV_X32 U_g13323 ( .A(I20390), .ZN(g13323) );
INV_X32 U_g13324 ( .A(g10316), .ZN(g13324) );
INV_X32 U_I20394 ( .A(g10331), .ZN(I20394) );
INV_X32 U_g13325 ( .A(I20394), .ZN(g13325) );
INV_X32 U_I20398 ( .A(g10858), .ZN(I20398) );
INV_X32 U_g13327 ( .A(I20398), .ZN(g13327) );
INV_X32 U_g13328 ( .A(g10334), .ZN(g13328) );
INV_X32 U_g13329 ( .A(g10337), .ZN(g13329) );
INV_X32 U_g13330 ( .A(g10357), .ZN(g13330) );
INV_X32 U_I20407 ( .A(g9027), .ZN(I20407) );
INV_X32 U_g13336 ( .A(I20407), .ZN(g13336) );
INV_X32 U_I20410 ( .A(g10887), .ZN(I20410) );
INV_X32 U_g13339 ( .A(I20410), .ZN(g13339) );
INV_X32 U_I20414 ( .A(g8575), .ZN(I20414) );
INV_X32 U_g13341 ( .A(I20414), .ZN(g13341) );
INV_X32 U_I20417 ( .A(g10933), .ZN(I20417) );
INV_X32 U_g13342 ( .A(I20417), .ZN(g13342) );
INV_X32 U_I20421 ( .A(g10808), .ZN(I20421) );
INV_X32 U_g13344 ( .A(I20421), .ZN(g13344) );
INV_X32 U_I20425 ( .A(g10842), .ZN(I20425) );
INV_X32 U_g13346 ( .A(I20425), .ZN(g13346) );
INV_X32 U_g13347 ( .A(g10409), .ZN(g13347) );
INV_X32 U_g13351 ( .A(g10416), .ZN(g13351) );
INV_X32 U_g13352 ( .A(g10419), .ZN(g13352) );
INV_X32 U_I20441 ( .A(g9027), .ZN(I20441) );
INV_X32 U_g13356 ( .A(I20441), .ZN(g13356) );
INV_X32 U_I20444 ( .A(g10869), .ZN(I20444) );
INV_X32 U_g13359 ( .A(I20444), .ZN(g13359) );
INV_X32 U_I20448 ( .A(g9050), .ZN(I20448) );
INV_X32 U_g13361 ( .A(I20448), .ZN(g13361) );
INV_X32 U_I20451 ( .A(g10908), .ZN(I20451) );
INV_X32 U_g13364 ( .A(I20451), .ZN(g13364) );
INV_X32 U_I20455 ( .A(g8578), .ZN(I20455) );
INV_X32 U_g13366 ( .A(I20455), .ZN(g13366) );
INV_X32 U_I20458 ( .A(g10972), .ZN(I20458) );
INV_X32 U_g13367 ( .A(I20458), .ZN(g13367) );
INV_X32 U_I20462 ( .A(g10825), .ZN(I20462) );
INV_X32 U_g13369 ( .A(I20462), .ZN(g13369) );
INV_X32 U_g13373 ( .A(g10482), .ZN(g13373) );
INV_X32 U_I20476 ( .A(g9027), .ZN(I20476) );
INV_X32 U_g13381 ( .A(I20476), .ZN(g13381) );
INV_X32 U_I20479 ( .A(g10849), .ZN(I20479) );
INV_X32 U_g13384 ( .A(I20479), .ZN(g13384) );
INV_X32 U_I20483 ( .A(g9050), .ZN(I20483) );
INV_X32 U_g13386 ( .A(I20483), .ZN(g13386) );
INV_X32 U_I20486 ( .A(g10889), .ZN(I20486) );
INV_X32 U_g13389 ( .A(I20486), .ZN(g13389) );
INV_X32 U_I20490 ( .A(g9067), .ZN(I20490) );
INV_X32 U_g13391 ( .A(I20490), .ZN(g13391) );
INV_X32 U_I20493 ( .A(g10934), .ZN(I20493) );
INV_X32 U_g13394 ( .A(I20493), .ZN(g13394) );
INV_X32 U_I20497 ( .A(g8579), .ZN(I20497) );
INV_X32 U_g13396 ( .A(I20497), .ZN(g13396) );
INV_X32 U_I20500 ( .A(g11007), .ZN(I20500) );
INV_X32 U_g13397 ( .A(I20500), .ZN(g13397) );
INV_X32 U_g13398 ( .A(g10542), .ZN(g13398) );
INV_X32 U_g13400 ( .A(g10545), .ZN(g13400) );
INV_X32 U_I20514 ( .A(g11769), .ZN(I20514) );
INV_X32 U_g13405 ( .A(I20514), .ZN(g13405) );
INV_X32 U_I20517 ( .A(g12425), .ZN(I20517) );
INV_X32 U_g13406 ( .A(I20517), .ZN(g13406) );
INV_X32 U_I20520 ( .A(g13246), .ZN(I20520) );
INV_X32 U_g13407 ( .A(I20520), .ZN(g13407) );
INV_X32 U_I20523 ( .A(g13317), .ZN(I20523) );
INV_X32 U_g13408 ( .A(I20523), .ZN(g13408) );
INV_X32 U_I20526 ( .A(g12519), .ZN(I20526) );
INV_X32 U_g13409 ( .A(I20526), .ZN(g13409) );
INV_X32 U_I20529 ( .A(g13319), .ZN(I20529) );
INV_X32 U_g13410 ( .A(I20529), .ZN(g13410) );
INV_X32 U_I20532 ( .A(g13339), .ZN(I20532) );
INV_X32 U_g13411 ( .A(I20532), .ZN(g13411) );
INV_X32 U_I20535 ( .A(g13359), .ZN(I20535) );
INV_X32 U_g13412 ( .A(I20535), .ZN(g13412) );
INV_X32 U_I20538 ( .A(g13384), .ZN(I20538) );
INV_X32 U_g13413 ( .A(I20538), .ZN(g13413) );
INV_X32 U_I20541 ( .A(g11599), .ZN(I20541) );
INV_X32 U_g13414 ( .A(I20541), .ZN(g13414) );
INV_X32 U_I20544 ( .A(g11628), .ZN(I20544) );
INV_X32 U_g13415 ( .A(I20544), .ZN(g13415) );
INV_X32 U_I20547 ( .A(g13248), .ZN(I20547) );
INV_X32 U_g13416 ( .A(I20547), .ZN(g13416) );
INV_X32 U_I20550 ( .A(g13267), .ZN(I20550) );
INV_X32 U_g13417 ( .A(I20550), .ZN(g13417) );
INV_X32 U_I20553 ( .A(g13290), .ZN(I20553) );
INV_X32 U_g13418 ( .A(I20553), .ZN(g13418) );
INV_X32 U_I20556 ( .A(g12435), .ZN(I20556) );
INV_X32 U_g13419 ( .A(I20556), .ZN(g13419) );
INV_X32 U_I20559 ( .A(g11937), .ZN(I20559) );
INV_X32 U_g13420 ( .A(I20559), .ZN(g13420) );
INV_X32 U_I20562 ( .A(g11786), .ZN(I20562) );
INV_X32 U_g13421 ( .A(I20562), .ZN(g13421) );
INV_X32 U_I20565 ( .A(g12432), .ZN(I20565) );
INV_X32 U_g13422 ( .A(I20565), .ZN(g13422) );
INV_X32 U_I20568 ( .A(g13269), .ZN(I20568) );
INV_X32 U_g13423 ( .A(I20568), .ZN(g13423) );
INV_X32 U_I20571 ( .A(g13341), .ZN(I20571) );
INV_X32 U_g13424 ( .A(I20571), .ZN(g13424) );
INV_X32 U_I20574 ( .A(g12534), .ZN(I20574) );
INV_X32 U_g13425 ( .A(I20574), .ZN(g13425) );
INV_X32 U_I20577 ( .A(g13342), .ZN(I20577) );
INV_X32 U_g13426 ( .A(I20577), .ZN(g13426) );
INV_X32 U_I20580 ( .A(g13364), .ZN(I20580) );
INV_X32 U_g13427 ( .A(I20580), .ZN(g13427) );
INV_X32 U_I20583 ( .A(g13389), .ZN(I20583) );
INV_X32 U_g13428 ( .A(I20583), .ZN(g13428) );
INV_X32 U_I20586 ( .A(g11606), .ZN(I20586) );
INV_X32 U_g13429 ( .A(I20586), .ZN(g13429) );
INV_X32 U_I20589 ( .A(g11629), .ZN(I20589) );
INV_X32 U_g13430 ( .A(I20589), .ZN(g13430) );
INV_X32 U_I20592 ( .A(g11651), .ZN(I20592) );
INV_X32 U_g13431 ( .A(I20592), .ZN(g13431) );
INV_X32 U_I20595 ( .A(g13271), .ZN(I20595) );
INV_X32 U_g13432 ( .A(I20595), .ZN(g13432) );
INV_X32 U_I20598 ( .A(g13292), .ZN(I20598) );
INV_X32 U_g13433 ( .A(I20598), .ZN(g13433) );
INV_X32 U_I20601 ( .A(g13321), .ZN(I20601) );
INV_X32 U_g13434 ( .A(I20601), .ZN(g13434) );
INV_X32 U_I20604 ( .A(g12440), .ZN(I20604) );
INV_X32 U_g13435 ( .A(I20604), .ZN(g13435) );
INV_X32 U_I20607 ( .A(g11990), .ZN(I20607) );
INV_X32 U_g13436 ( .A(I20607), .ZN(g13436) );
INV_X32 U_I20610 ( .A(g11812), .ZN(I20610) );
INV_X32 U_g13437 ( .A(I20610), .ZN(g13437) );
INV_X32 U_I20613 ( .A(g12437), .ZN(I20613) );
INV_X32 U_g13438 ( .A(I20613), .ZN(g13438) );
INV_X32 U_I20616 ( .A(g13294), .ZN(I20616) );
INV_X32 U_g13439 ( .A(I20616), .ZN(g13439) );
INV_X32 U_I20619 ( .A(g13366), .ZN(I20619) );
INV_X32 U_g13440 ( .A(I20619), .ZN(g13440) );
INV_X32 U_I20622 ( .A(g12543), .ZN(I20622) );
INV_X32 U_g13441 ( .A(I20622), .ZN(g13441) );
INV_X32 U_I20625 ( .A(g13367), .ZN(I20625) );
INV_X32 U_g13442 ( .A(I20625), .ZN(g13442) );
INV_X32 U_I20628 ( .A(g13394), .ZN(I20628) );
INV_X32 U_g13443 ( .A(I20628), .ZN(g13443) );
INV_X32 U_I20631 ( .A(g11611), .ZN(I20631) );
INV_X32 U_g13444 ( .A(I20631), .ZN(g13444) );
INV_X32 U_I20634 ( .A(g11636), .ZN(I20634) );
INV_X32 U_g13445 ( .A(I20634), .ZN(g13445) );
INV_X32 U_I20637 ( .A(g11652), .ZN(I20637) );
INV_X32 U_g13446 ( .A(I20637), .ZN(g13446) );
INV_X32 U_I20640 ( .A(g11670), .ZN(I20640) );
INV_X32 U_g13447 ( .A(I20640), .ZN(g13447) );
INV_X32 U_I20643 ( .A(g13296), .ZN(I20643) );
INV_X32 U_g13448 ( .A(I20643), .ZN(g13448) );
INV_X32 U_I20646 ( .A(g13323), .ZN(I20646) );
INV_X32 U_g13449 ( .A(I20646), .ZN(g13449) );
INV_X32 U_I20649 ( .A(g13344), .ZN(I20649) );
INV_X32 U_g13450 ( .A(I20649), .ZN(g13450) );
INV_X32 U_I20652 ( .A(g12445), .ZN(I20652) );
INV_X32 U_g13451 ( .A(I20652), .ZN(g13451) );
INV_X32 U_I20655 ( .A(g12059), .ZN(I20655) );
INV_X32 U_g13452 ( .A(I20655), .ZN(g13452) );
INV_X32 U_I20658 ( .A(g11845), .ZN(I20658) );
INV_X32 U_g13453 ( .A(I20658), .ZN(g13453) );
INV_X32 U_I20661 ( .A(g12442), .ZN(I20661) );
INV_X32 U_g13454 ( .A(I20661), .ZN(g13454) );
INV_X32 U_I20664 ( .A(g13325), .ZN(I20664) );
INV_X32 U_g13455 ( .A(I20664), .ZN(g13455) );
INV_X32 U_I20667 ( .A(g13396), .ZN(I20667) );
INV_X32 U_g13456 ( .A(I20667), .ZN(g13456) );
INV_X32 U_I20670 ( .A(g12552), .ZN(I20670) );
INV_X32 U_g13457 ( .A(I20670), .ZN(g13457) );
INV_X32 U_I20673 ( .A(g13397), .ZN(I20673) );
INV_X32 U_g13458 ( .A(I20673), .ZN(g13458) );
INV_X32 U_I20676 ( .A(g11616), .ZN(I20676) );
INV_X32 U_g13459 ( .A(I20676), .ZN(g13459) );
INV_X32 U_I20679 ( .A(g11641), .ZN(I20679) );
INV_X32 U_g13460 ( .A(I20679), .ZN(g13460) );
INV_X32 U_I20682 ( .A(g11659), .ZN(I20682) );
INV_X32 U_g13461 ( .A(I20682), .ZN(g13461) );
INV_X32 U_I20685 ( .A(g11671), .ZN(I20685) );
INV_X32 U_g13462 ( .A(I20685), .ZN(g13462) );
INV_X32 U_I20688 ( .A(g11682), .ZN(I20688) );
INV_X32 U_g13463 ( .A(I20688), .ZN(g13463) );
INV_X32 U_I20691 ( .A(g13327), .ZN(I20691) );
INV_X32 U_g13464 ( .A(I20691), .ZN(g13464) );
INV_X32 U_I20694 ( .A(g13346), .ZN(I20694) );
INV_X32 U_g13465 ( .A(I20694), .ZN(g13465) );
INV_X32 U_I20697 ( .A(g13369), .ZN(I20697) );
INV_X32 U_g13466 ( .A(I20697), .ZN(g13466) );
INV_X32 U_I20700 ( .A(g12450), .ZN(I20700) );
INV_X32 U_g13467 ( .A(I20700), .ZN(g13467) );
INV_X32 U_I20703 ( .A(g12123), .ZN(I20703) );
INV_X32 U_g13468 ( .A(I20703), .ZN(g13468) );
INV_X32 U_I20706 ( .A(g11490), .ZN(I20706) );
INV_X32 U_g13469 ( .A(I20706), .ZN(g13469) );
INV_X32 U_I20709 ( .A(g13070), .ZN(I20709) );
INV_X32 U_g13475 ( .A(I20709), .ZN(g13475) );
INV_X32 U_g13519 ( .A(g13228), .ZN(g13519) );
INV_X32 U_g13530 ( .A(g13251), .ZN(g13530) );
INV_X32 U_g13541 ( .A(g13274), .ZN(g13541) );
INV_X32 U_g13552 ( .A(g13299), .ZN(g13552) );
INV_X32 U_g13565 ( .A(g12192), .ZN(g13565) );
INV_X32 U_g13568 ( .A(g11627), .ZN(g13568) );
INV_X32 U_I20791 ( .A(g13149), .ZN(I20791) );
INV_X32 U_g13571 ( .A(I20791), .ZN(g13571) );
INV_X32 U_I20794 ( .A(g13111), .ZN(I20794) );
INV_X32 U_g13572 ( .A(I20794), .ZN(g13572) );
INV_X32 U_g13573 ( .A(g12247), .ZN(g13573) );
INV_X32 U_g13576 ( .A(g11650), .ZN(g13576) );
INV_X32 U_I20799 ( .A(g13155), .ZN(I20799) );
INV_X32 U_g13579 ( .A(I20799), .ZN(g13579) );
INV_X32 U_I20802 ( .A(g13160), .ZN(I20802) );
INV_X32 U_g13580 ( .A(I20802), .ZN(g13580) );
INV_X32 U_I20805 ( .A(g13124), .ZN(I20805) );
INV_X32 U_g13581 ( .A(I20805), .ZN(g13581) );
INV_X32 U_g13582 ( .A(g12290), .ZN(g13582) );
INV_X32 U_g13585 ( .A(g11669), .ZN(g13585) );
INV_X32 U_I20810 ( .A(g13164), .ZN(I20810) );
INV_X32 U_g13588 ( .A(I20810), .ZN(g13588) );
INV_X32 U_I20813 ( .A(g13265), .ZN(I20813) );
INV_X32 U_g13589 ( .A(I20813), .ZN(g13589) );
INV_X32 U_I20816 ( .A(g12487), .ZN(I20816) );
INV_X32 U_g13598 ( .A(I20816), .ZN(g13598) );
INV_X32 U_I20820 ( .A(g13171), .ZN(I20820) );
INV_X32 U_g13600 ( .A(I20820), .ZN(g13600) );
INV_X32 U_I20823 ( .A(g13135), .ZN(I20823) );
INV_X32 U_g13601 ( .A(I20823), .ZN(g13601) );
INV_X32 U_g13602 ( .A(g12326), .ZN(g13602) );
INV_X32 U_g13605 ( .A(g11681), .ZN(g13605) );
INV_X32 U_I20828 ( .A(g13175), .ZN(I20828) );
INV_X32 U_g13608 ( .A(I20828), .ZN(g13608) );
INV_X32 U_I20832 ( .A(g12507), .ZN(I20832) );
INV_X32 U_g13610 ( .A(I20832), .ZN(g13610) );
INV_X32 U_I20836 ( .A(g13182), .ZN(I20836) );
INV_X32 U_g13612 ( .A(I20836), .ZN(g13612) );
INV_X32 U_I20839 ( .A(g13143), .ZN(I20839) );
INV_X32 U_g13613 ( .A(I20839), .ZN(g13613) );
INV_X32 U_g13614 ( .A(g11690), .ZN(g13614) );
INV_X32 U_I20844 ( .A(g12524), .ZN(I20844) );
INV_X32 U_g13620 ( .A(I20844), .ZN(g13620) );
INV_X32 U_I20848 ( .A(g13194), .ZN(I20848) );
INV_X32 U_g13622 ( .A(I20848), .ZN(g13622) );
INV_X32 U_I20852 ( .A(g12457), .ZN(I20852) );
INV_X32 U_g13624 ( .A(I20852), .ZN(g13624) );
INV_X32 U_g13626 ( .A(g11697), .ZN(g13626) );
INV_X32 U_I20858 ( .A(g12539), .ZN(I20858) );
INV_X32 U_g13632 ( .A(I20858), .ZN(g13632) );
INV_X32 U_I20863 ( .A(g12467), .ZN(I20863) );
INV_X32 U_g13635 ( .A(I20863), .ZN(g13635) );
INV_X32 U_g13637 ( .A(g11703), .ZN(g13637) );
INV_X32 U_g13644 ( .A(g13215), .ZN(g13644) );
INV_X32 U_I20873 ( .A(g12482), .ZN(I20873) );
INV_X32 U_g13647 ( .A(I20873), .ZN(g13647) );
INV_X32 U_g13649 ( .A(g11711), .ZN(g13649) );
INV_X32 U_g13657 ( .A(g12452), .ZN(g13657) );
INV_X32 U_g13669 ( .A(g13229), .ZN(g13669) );
INV_X32 U_g13670 ( .A(g13234), .ZN(g13670) );
INV_X32 U_I20886 ( .A(g12499), .ZN(I20886) );
INV_X32 U_g13673 ( .A(I20886), .ZN(g13673) );
INV_X32 U_g13677 ( .A(g12447), .ZN(g13677) );
INV_X32 U_g13687 ( .A(g12460), .ZN(g13687) );
INV_X32 U_g13699 ( .A(g13252), .ZN(g13699) );
INV_X32 U_g13700 ( .A(g13257), .ZN(g13700) );
INV_X32 U_g13706 ( .A(g12443), .ZN(g13706) );
INV_X32 U_g13714 ( .A(g12453), .ZN(g13714) );
INV_X32 U_g13724 ( .A(g12470), .ZN(g13724) );
INV_X32 U_g13736 ( .A(g13275), .ZN(g13736) );
INV_X32 U_g13737 ( .A(g13280), .ZN(g13737) );
INV_X32 U_I20909 ( .A(g13055), .ZN(I20909) );
INV_X32 U_g13741 ( .A(I20909), .ZN(g13741) );
INV_X32 U_g13750 ( .A(g12439), .ZN(g13750) );
INV_X32 U_g13756 ( .A(g12448), .ZN(g13756) );
INV_X32 U_g13764 ( .A(g12461), .ZN(g13764) );
INV_X32 U_g13774 ( .A(g12485), .ZN(g13774) );
INV_X32 U_g13786 ( .A(g13300), .ZN(g13786) );
INV_X32 U_g13791 ( .A(g12444), .ZN(g13791) );
INV_X32 U_g13797 ( .A(g12454), .ZN(g13797) );
INV_X32 U_g13805 ( .A(g12471), .ZN(g13805) );
INV_X32 U_g13817 ( .A(g13336), .ZN(g13817) );
INV_X32 U_g13819 ( .A(g12449), .ZN(g13819) );
INV_X32 U_g13825 ( .A(g12462), .ZN(g13825) );
INV_X32 U_g13836 ( .A(g13356), .ZN(g13836) );
INV_X32 U_g13838 ( .A(g13361), .ZN(g13838) );
INV_X32 U_g13840 ( .A(g12455), .ZN(g13840) );
INV_X32 U_g13848 ( .A(g11744), .ZN(g13848) );
INV_X32 U_g13849 ( .A(g13381), .ZN(g13849) );
INV_X32 U_g13850 ( .A(g13386), .ZN(g13850) );
INV_X32 U_g13852 ( .A(g13391), .ZN(g13852) );
INV_X32 U_g13856 ( .A(g11759), .ZN(g13856) );
INV_X32 U_g13857 ( .A(g11760), .ZN(g13857) );
INV_X32 U_g13858 ( .A(g11603), .ZN(g13858) );
INV_X32 U_g13859 ( .A(g11608), .ZN(g13859) );
INV_X32 U_g13861 ( .A(g11613), .ZN(g13861) );
INV_X32 U_I20959 ( .A(g11713), .ZN(I20959) );
INV_X32 U_g13863 ( .A(I20959), .ZN(g13863) );
INV_X32 U_g13864 ( .A(g11767), .ZN(g13864) );
INV_X32 U_g13866 ( .A(g11772), .ZN(g13866) );
INV_X32 U_g13867 ( .A(g11773), .ZN(g13867) );
INV_X32 U_g13868 ( .A(g11633), .ZN(g13868) );
INV_X32 U_g13869 ( .A(g11638), .ZN(g13869) );
INV_X32 U_g13872 ( .A(g11780), .ZN(g13872) );
INV_X32 U_g13873 ( .A(g12698), .ZN(g13873) );
INV_X32 U_g13879 ( .A(g11784), .ZN(g13879) );
INV_X32 U_g13881 ( .A(g11789), .ZN(g13881) );
INV_X32 U_g13882 ( .A(g11790), .ZN(g13882) );
INV_X32 U_g13883 ( .A(g11656), .ZN(g13883) );
INV_X32 U_g13885 ( .A(g11799), .ZN(g13885) );
INV_X32 U_g13886 ( .A(g12747), .ZN(g13886) );
INV_X32 U_g13894 ( .A(g11806), .ZN(g13894) );
INV_X32 U_g13895 ( .A(g12755), .ZN(g13895) );
INV_X32 U_g13901 ( .A(g11810), .ZN(g13901) );
INV_X32 U_g13903 ( .A(g11815), .ZN(g13903) );
INV_X32 U_g13906 ( .A(g11822), .ZN(g13906) );
INV_X32 U_g13907 ( .A(g12781), .ZN(g13907) );
INV_X32 U_g13918 ( .A(g11830), .ZN(g13918) );
INV_X32 U_g13922 ( .A(g11831), .ZN(g13922) );
INV_X32 U_g13926 ( .A(g11832), .ZN(g13926) );
INV_X32 U_g13927 ( .A(g12789), .ZN(g13927) );
INV_X32 U_g13935 ( .A(g11839), .ZN(g13935) );
INV_X32 U_g13936 ( .A(g12797), .ZN(g13936) );
INV_X32 U_g13942 ( .A(g11843), .ZN(g13942) );
INV_X32 U_g13945 ( .A(g11855), .ZN(g13945) );
INV_X32 U_g13946 ( .A(g12814), .ZN(g13946) );
INV_X32 U_I21012 ( .A(g12503), .ZN(I21012) );
INV_X32 U_g13954 ( .A(I21012), .ZN(g13954) );
INV_X32 U_g13958 ( .A(g11863), .ZN(g13958) );
INV_X32 U_g13962 ( .A(g11864), .ZN(g13962) );
INV_X32 U_g13963 ( .A(g12820), .ZN(g13963) );
INV_X32 U_g13974 ( .A(g11872), .ZN(g13974) );
INV_X32 U_g13978 ( .A(g11873), .ZN(g13978) );
INV_X32 U_g13982 ( .A(g11874), .ZN(g13982) );
INV_X32 U_g13983 ( .A(g12828), .ZN(g13983) );
INV_X32 U_g13991 ( .A(g11881), .ZN(g13991) );
INV_X32 U_g13992 ( .A(g12836), .ZN(g13992) );
INV_X32 U_g13999 ( .A(g11889), .ZN(g13999) );
INV_X32 U_g14000 ( .A(g11890), .ZN(g14000) );
INV_X32 U_g14001 ( .A(g12849), .ZN(g14001) );
INV_X32 U_I21037 ( .A(g12486), .ZN(I21037) );
INV_X32 U_g14008 ( .A(I21037), .ZN(g14008) );
INV_X32 U_g14011 ( .A(g11896), .ZN(g14011) );
INV_X32 U_g14015 ( .A(g11897), .ZN(g14015) );
INV_X32 U_g14016 ( .A(g12852), .ZN(g14016) );
INV_X32 U_I21045 ( .A(g12520), .ZN(I21045) );
INV_X32 U_g14024 ( .A(I21045), .ZN(g14024) );
INV_X32 U_g14028 ( .A(g11905), .ZN(g14028) );
INV_X32 U_g14032 ( .A(g11906), .ZN(g14032) );
INV_X32 U_g14033 ( .A(g12858), .ZN(g14033) );
INV_X32 U_g14044 ( .A(g11914), .ZN(g14044) );
INV_X32 U_g14048 ( .A(g11915), .ZN(g14048) );
INV_X32 U_g14052 ( .A(g11916), .ZN(g14052) );
INV_X32 U_g14053 ( .A(g12866), .ZN(g14053) );
INV_X32 U_g14061 ( .A(g11928), .ZN(g14061) );
INV_X32 U_g14062 ( .A(g12880), .ZN(g14062) );
INV_X32 U_I21064 ( .A(g13147), .ZN(I21064) );
INV_X32 U_g14068 ( .A(I21064), .ZN(g14068) );
INV_X32 U_g14071 ( .A(g11934), .ZN(g14071) );
INV_X32 U_g14079 ( .A(g11935), .ZN(g14079) );
INV_X32 U_g14086 ( .A(g11938), .ZN(g14086) );
INV_X32 U_g14090 ( .A(g11939), .ZN(g14090) );
INV_X32 U_g14091 ( .A(g11940), .ZN(g14091) );
INV_X32 U_g14092 ( .A(g12890), .ZN(g14092) );
INV_X32 U_I21075 ( .A(g12506), .ZN(I21075) );
INV_X32 U_g14099 ( .A(I21075), .ZN(g14099) );
INV_X32 U_g14102 ( .A(g11946), .ZN(g14102) );
INV_X32 U_g14106 ( .A(g11947), .ZN(g14106) );
INV_X32 U_g14107 ( .A(g12893), .ZN(g14107) );
INV_X32 U_I21083 ( .A(g12535), .ZN(I21083) );
INV_X32 U_g14115 ( .A(I21083), .ZN(g14115) );
INV_X32 U_g14119 ( .A(g11955), .ZN(g14119) );
INV_X32 U_g14123 ( .A(g11956), .ZN(g14123) );
INV_X32 U_g14124 ( .A(g12899), .ZN(g14124) );
INV_X32 U_g14135 ( .A(g11964), .ZN(g14135) );
INV_X32 U_g14139 ( .A(g11965), .ZN(g14139) );
INV_X32 U_I21096 ( .A(g11749), .ZN(I21096) );
INV_X32 U_g14144 ( .A(I21096), .ZN(g14144) );
INV_X32 U_g14148 ( .A(g12912), .ZN(g14148) );
INV_X32 U_g14153 ( .A(g12913), .ZN(g14153) );
INV_X32 U_g14158 ( .A(g11974), .ZN(g14158) );
INV_X32 U_g14165 ( .A(g11975), .ZN(g14165) );
INV_X32 U_g14171 ( .A(g11979), .ZN(g14171) );
INV_X32 U_g14175 ( .A(g11980), .ZN(g14175) );
INV_X32 U_g14176 ( .A(g11981), .ZN(g14176) );
INV_X32 U_g14177 ( .A(g12920), .ZN(g14177) );
INV_X32 U_I21108 ( .A(g13150), .ZN(I21108) );
INV_X32 U_g14183 ( .A(I21108), .ZN(g14183) );
INV_X32 U_g14186 ( .A(g11987), .ZN(g14186) );
INV_X32 U_g14194 ( .A(g11988), .ZN(g14194) );
INV_X32 U_g14201 ( .A(g11991), .ZN(g14201) );
INV_X32 U_g14205 ( .A(g11992), .ZN(g14205) );
INV_X32 U_g14206 ( .A(g11993), .ZN(g14206) );
INV_X32 U_g14207 ( .A(g12930), .ZN(g14207) );
INV_X32 U_I21119 ( .A(g12523), .ZN(I21119) );
INV_X32 U_g14214 ( .A(I21119), .ZN(g14214) );
INV_X32 U_g14217 ( .A(g11999), .ZN(g14217) );
INV_X32 U_g14221 ( .A(g12000), .ZN(g14221) );
INV_X32 U_g14222 ( .A(g12933), .ZN(g14222) );
INV_X32 U_I21127 ( .A(g12544), .ZN(I21127) );
INV_X32 U_g14230 ( .A(I21127), .ZN(g14230) );
INV_X32 U_g14234 ( .A(g12008), .ZN(g14234) );
INV_X32 U_g14238 ( .A(g12939), .ZN(g14238) );
INV_X32 U_g14244 ( .A(g12026), .ZN(g14244) );
INV_X32 U_g14249 ( .A(g12034), .ZN(g14249) );
INV_X32 U_g14252 ( .A(g12035), .ZN(g14252) );
INV_X32 U_g14256 ( .A(g12036), .ZN(g14256) );
INV_X32 U_I21137 ( .A(g11749), .ZN(I21137) );
INV_X32 U_g14259 ( .A(I21137), .ZN(g14259) );
INV_X32 U_g14263 ( .A(g12941), .ZN(g14263) );
INV_X32 U_g14268 ( .A(g12942), .ZN(g14268) );
INV_X32 U_g14273 ( .A(g12043), .ZN(g14273) );
INV_X32 U_g14280 ( .A(g12044), .ZN(g14280) );
INV_X32 U_g14286 ( .A(g12048), .ZN(g14286) );
INV_X32 U_g14290 ( .A(g12049), .ZN(g14290) );
INV_X32 U_g14291 ( .A(g12050), .ZN(g14291) );
INV_X32 U_g14292 ( .A(g12949), .ZN(g14292) );
INV_X32 U_I21149 ( .A(g13156), .ZN(I21149) );
INV_X32 U_g14298 ( .A(I21149), .ZN(g14298) );
INV_X32 U_g14301 ( .A(g12056), .ZN(g14301) );
INV_X32 U_g14309 ( .A(g12057), .ZN(g14309) );
INV_X32 U_g14316 ( .A(g12060), .ZN(g14316) );
INV_X32 U_g14320 ( .A(g12061), .ZN(g14320) );
INV_X32 U_g14321 ( .A(g12062), .ZN(g14321) );
INV_X32 U_g14322 ( .A(g12959), .ZN(g14322) );
INV_X32 U_I21160 ( .A(g12538), .ZN(I21160) );
INV_X32 U_g14329 ( .A(I21160), .ZN(g14329) );
INV_X32 U_g14332 ( .A(g12068), .ZN(g14332) );
INV_X32 U_I21165 ( .A(g13110), .ZN(I21165) );
INV_X32 U_g14337 ( .A(I21165), .ZN(g14337) );
INV_X32 U_g14342 ( .A(g12967), .ZN(g14342) );
INV_X32 U_g14347 ( .A(g12079), .ZN(g14347) );
INV_X32 U_g14352 ( .A(g12081), .ZN(g14352) );
INV_X32 U_g14355 ( .A(g12082), .ZN(g14355) );
INV_X32 U_g14359 ( .A(g12083), .ZN(g14359) );
INV_X32 U_g14360 ( .A(g12968), .ZN(g14360) );
INV_X32 U_g14366 ( .A(g12090), .ZN(g14366) );
INV_X32 U_g14371 ( .A(g12098), .ZN(g14371) );
INV_X32 U_g14374 ( .A(g12099), .ZN(g14374) );
INV_X32 U_g14378 ( .A(g12100), .ZN(g14378) );
INV_X32 U_I21178 ( .A(g11749), .ZN(I21178) );
INV_X32 U_g14381 ( .A(I21178), .ZN(g14381) );
INV_X32 U_g14385 ( .A(g12970), .ZN(g14385) );
INV_X32 U_g14390 ( .A(g12971), .ZN(g14390) );
INV_X32 U_g14395 ( .A(g12107), .ZN(g14395) );
INV_X32 U_g14402 ( .A(g12108), .ZN(g14402) );
INV_X32 U_g14408 ( .A(g12112), .ZN(g14408) );
INV_X32 U_g14412 ( .A(g12113), .ZN(g14412) );
INV_X32 U_g14413 ( .A(g12114), .ZN(g14413) );
INV_X32 U_g14414 ( .A(g12978), .ZN(g14414) );
INV_X32 U_I21190 ( .A(g13165), .ZN(I21190) );
INV_X32 U_g14420 ( .A(I21190), .ZN(g14420) );
INV_X32 U_g14423 ( .A(g12120), .ZN(g14423) );
INV_X32 U_g14431 ( .A(g12121), .ZN(g14431) );
INV_X32 U_g14438 ( .A(g12124), .ZN(g14438) );
INV_X32 U_g14442 ( .A(g11768), .ZN(g14442) );
INV_X32 U_g14450 ( .A(g12146), .ZN(g14450) );
INV_X32 U_g14454 ( .A(g12991), .ZN(g14454) );
INV_X32 U_g14459 ( .A(g12151), .ZN(g14459) );
INV_X32 U_g14464 ( .A(g12153), .ZN(g14464) );
INV_X32 U_g14467 ( .A(g12154), .ZN(g14467) );
INV_X32 U_g14471 ( .A(g12155), .ZN(g14471) );
INV_X32 U_g14472 ( .A(g12992), .ZN(g14472) );
INV_X32 U_g14478 ( .A(g12162), .ZN(g14478) );
INV_X32 U_g14483 ( .A(g12170), .ZN(g14483) );
INV_X32 U_g14486 ( .A(g12171), .ZN(g14486) );
INV_X32 U_g14490 ( .A(g12172), .ZN(g14490) );
INV_X32 U_I21208 ( .A(g11749), .ZN(I21208) );
INV_X32 U_g14493 ( .A(I21208), .ZN(g14493) );
INV_X32 U_g14497 ( .A(g12994), .ZN(g14497) );
INV_X32 U_g14502 ( .A(g12995), .ZN(g14502) );
INV_X32 U_g14507 ( .A(g12179), .ZN(g14507) );
INV_X32 U_g14514 ( .A(g12180), .ZN(g14514) );
INV_X32 U_g14520 ( .A(g12184), .ZN(g14520) );
INV_X32 U_g14524 ( .A(g12185), .ZN(g14524) );
INV_X32 U_g14525 ( .A(g12195), .ZN(g14525) );
INV_X32 U_g14529 ( .A(g11785), .ZN(g14529) );
INV_X32 U_g14537 ( .A(g12208), .ZN(g14537) );
INV_X32 U_g14541 ( .A(g13001), .ZN(g14541) );
INV_X32 U_g14546 ( .A(g12213), .ZN(g14546) );
INV_X32 U_g14551 ( .A(g12215), .ZN(g14551) );
INV_X32 U_g14554 ( .A(g12216), .ZN(g14554) );
INV_X32 U_g14558 ( .A(g12217), .ZN(g14558) );
INV_X32 U_g14559 ( .A(g13002), .ZN(g14559) );
INV_X32 U_g14565 ( .A(g12224), .ZN(g14565) );
INV_X32 U_g14570 ( .A(g12232), .ZN(g14570) );
INV_X32 U_g14573 ( .A(g12233), .ZN(g14573) );
INV_X32 U_g14577 ( .A(g12234), .ZN(g14577) );
INV_X32 U_g14580 ( .A(g12250), .ZN(g14580) );
INV_X32 U_g14584 ( .A(g11811), .ZN(g14584) );
INV_X32 U_g14592 ( .A(g12263), .ZN(g14592) );
INV_X32 U_g14596 ( .A(g13022), .ZN(g14596) );
INV_X32 U_g14601 ( .A(g12268), .ZN(g14601) );
INV_X32 U_g14606 ( .A(g12270), .ZN(g14606) );
INV_X32 U_g14609 ( .A(g12271), .ZN(g14609) );
INV_X32 U_g14613 ( .A(g12272), .ZN(g14613) );
INV_X32 U_g14614 ( .A(g12293), .ZN(g14614) );
INV_X32 U_g14618 ( .A(g11844), .ZN(g14618) );
INV_X32 U_g14626 ( .A(g12306), .ZN(g14626) );
INV_X32 U_I21241 ( .A(g13378), .ZN(I21241) );
INV_X32 U_g14630 ( .A(I21241), .ZN(g14630) );
INV_X32 U_g14637 ( .A(g12329), .ZN(g14637) );
INV_X32 U_g14641 ( .A(g11823), .ZN(g14641) );
INV_X32 U_I21246 ( .A(g11624), .ZN(I21246) );
INV_X32 U_g14642 ( .A(I21246), .ZN(g14642) );
INV_X32 U_I21249 ( .A(g11600), .ZN(I21249) );
INV_X32 U_g14650 ( .A(I21249), .ZN(g14650) );
INV_X32 U_I21252 ( .A(g11644), .ZN(I21252) );
INV_X32 U_g14657 ( .A(I21252), .ZN(g14657) );
INV_X32 U_g14668 ( .A(g11865), .ZN(g14668) );
INV_X32 U_I21256 ( .A(g11647), .ZN(I21256) );
INV_X32 U_g14669 ( .A(I21256), .ZN(g14669) );
INV_X32 U_I21259 ( .A(g11630), .ZN(I21259) );
INV_X32 U_g14677 ( .A(I21259), .ZN(g14677) );
INV_X32 U_I21262 ( .A(g11713), .ZN(I21262) );
INV_X32 U_g14684 ( .A(I21262), .ZN(g14684) );
INV_X32 U_g14685 ( .A(g12245), .ZN(g14685) );
INV_X32 U_I21267 ( .A(g11663), .ZN(I21267) );
INV_X32 U_g14691 ( .A(I21267), .ZN(g14691) );
INV_X32 U_g14702 ( .A(g11907), .ZN(g14702) );
INV_X32 U_I21271 ( .A(g11666), .ZN(I21271) );
INV_X32 U_g14703 ( .A(I21271), .ZN(g14703) );
INV_X32 U_I21274 ( .A(g11653), .ZN(I21274) );
INV_X32 U_g14711 ( .A(I21274), .ZN(g14711) );
INV_X32 U_I21277 ( .A(g12430), .ZN(I21277) );
INV_X32 U_g14718 ( .A(I21277), .ZN(g14718) );
INV_X32 U_g14719 ( .A(g12288), .ZN(g14719) );
INV_X32 U_I21282 ( .A(g11675), .ZN(I21282) );
INV_X32 U_g14725 ( .A(I21282), .ZN(g14725) );
INV_X32 U_g14736 ( .A(g11957), .ZN(g14736) );
INV_X32 U_I21286 ( .A(g11678), .ZN(I21286) );
INV_X32 U_g14737 ( .A(I21286), .ZN(g14737) );
INV_X32 U_I21289 ( .A(g12434), .ZN(I21289) );
INV_X32 U_g14745 ( .A(I21289), .ZN(g14745) );
INV_X32 U_I21292 ( .A(g11888), .ZN(I21292) );
INV_X32 U_g14746 ( .A(I21292), .ZN(g14746) );
INV_X32 U_g14747 ( .A(g12324), .ZN(g14747) );
INV_X32 U_I21297 ( .A(g11687), .ZN(I21297) );
INV_X32 U_g14753 ( .A(I21297), .ZN(g14753) );
INV_X32 U_g14764 ( .A(g11791), .ZN(g14764) );
INV_X32 U_I21301 ( .A(g12438), .ZN(I21301) );
INV_X32 U_g14765 ( .A(I21301), .ZN(g14765) );
INV_X32 U_I21304 ( .A(g11927), .ZN(I21304) );
INV_X32 U_g14766 ( .A(I21304), .ZN(g14766) );
INV_X32 U_g14768 ( .A(g12352), .ZN(g14768) );
INV_X32 U_I21310 ( .A(g12332), .ZN(I21310) );
INV_X32 U_g14774 ( .A(I21310), .ZN(g14774) );
INV_X32 U_I21313 ( .A(g11743), .ZN(I21313) );
INV_X32 U_g14775 ( .A(I21313), .ZN(g14775) );
INV_X32 U_g14776 ( .A(g12033), .ZN(g14776) );
INV_X32 U_g14794 ( .A(g11848), .ZN(g14794) );
INV_X32 U_I21318 ( .A(g12362), .ZN(I21318) );
INV_X32 U_g14795 ( .A(I21318), .ZN(g14795) );
INV_X32 U_I21321 ( .A(g11758), .ZN(I21321) );
INV_X32 U_g14796 ( .A(I21321), .ZN(g14796) );
INV_X32 U_g14797 ( .A(g12080), .ZN(g14797) );
INV_X32 U_g14811 ( .A(g12097), .ZN(g14811) );
INV_X32 U_I21326 ( .A(g12378), .ZN(I21326) );
INV_X32 U_g14829 ( .A(I21326), .ZN(g14829) );
INV_X32 U_I21329 ( .A(g11766), .ZN(I21329) );
INV_X32 U_g14830 ( .A(I21329), .ZN(g14830) );
INV_X32 U_g14831 ( .A(g11828), .ZN(g14831) );
INV_X32 U_g14837 ( .A(g12145), .ZN(g14837) );
INV_X32 U_g14849 ( .A(g12152), .ZN(g14849) );
INV_X32 U_g14863 ( .A(g12169), .ZN(g14863) );
INV_X32 U_g14881 ( .A(g11923), .ZN(g14881) );
INV_X32 U_I21337 ( .A(g12408), .ZN(I21337) );
INV_X32 U_g14882 ( .A(I21337), .ZN(g14882) );
INV_X32 U_I21340 ( .A(g11779), .ZN(I21340) );
INV_X32 U_g14883 ( .A(I21340), .ZN(g14883) );
INV_X32 U_g14885 ( .A(g11860), .ZN(g14885) );
INV_X32 U_g14895 ( .A(g12193), .ZN(g14895) );
INV_X32 U_g14904 ( .A(g11870), .ZN(g14904) );
INV_X32 U_g14910 ( .A(g12207), .ZN(g14910) );
INV_X32 U_g14922 ( .A(g12214), .ZN(g14922) );
INV_X32 U_g14936 ( .A(g12231), .ZN(g14936) );
INV_X32 U_I21351 ( .A(g12420), .ZN(I21351) );
INV_X32 U_g14954 ( .A(I21351), .ZN(g14954) );
INV_X32 U_I21354 ( .A(g11798), .ZN(I21354) );
INV_X32 U_g14955 ( .A(I21354), .ZN(g14955) );
INV_X32 U_g14959 ( .A(g11976), .ZN(g14959) );
INV_X32 U_I21361 ( .A(g13026), .ZN(I21361) );
INV_X32 U_g14960 ( .A(I21361), .ZN(g14960) );
INV_X32 U_I21364 ( .A(g13028), .ZN(I21364) );
INV_X32 U_g14963 ( .A(I21364), .ZN(g14963) );
INV_X32 U_g14966 ( .A(g11902), .ZN(g14966) );
INV_X32 U_g14976 ( .A(g12248), .ZN(g14976) );
INV_X32 U_g14985 ( .A(g11912), .ZN(g14985) );
INV_X32 U_g14991 ( .A(g12262), .ZN(g14991) );
INV_X32 U_g15003 ( .A(g12269), .ZN(g15003) );
INV_X32 U_g15017 ( .A(g12009), .ZN(g15017) );
INV_X32 U_I21374 ( .A(g12424), .ZN(I21374) );
INV_X32 U_g15018 ( .A(I21374), .ZN(g15018) );
INV_X32 U_I21377 ( .A(g11821), .ZN(I21377) );
INV_X32 U_g15019 ( .A(I21377), .ZN(g15019) );
INV_X32 U_I21381 ( .A(g13157), .ZN(I21381) );
INV_X32 U_g15021 ( .A(I21381), .ZN(g15021) );
INV_X32 U_g15022 ( .A(g11781), .ZN(g15022) );
INV_X32 U_g15032 ( .A(g12027), .ZN(g15032) );
INV_X32 U_g15033 ( .A(g12030), .ZN(g15033) );
INV_X32 U_I21389 ( .A(g12883), .ZN(I21389) );
INV_X32 U_g15034 ( .A(I21389), .ZN(g15034) );
INV_X32 U_I21392 ( .A(g13020), .ZN(I21392) );
INV_X32 U_g15037 ( .A(I21392), .ZN(g15037) );
INV_X32 U_I21395 ( .A(g13034), .ZN(I21395) );
INV_X32 U_g15040 ( .A(I21395), .ZN(g15040) );
INV_X32 U_I21398 ( .A(g13021), .ZN(I21398) );
INV_X32 U_g15043 ( .A(I21398), .ZN(g15043) );
INV_X32 U_g15048 ( .A(g12045), .ZN(g15048) );
INV_X32 U_I21404 ( .A(g13037), .ZN(I21404) );
INV_X32 U_g15049 ( .A(I21404), .ZN(g15049) );
INV_X32 U_I21407 ( .A(g13039), .ZN(I21407) );
INV_X32 U_g15052 ( .A(I21407), .ZN(g15052) );
INV_X32 U_g15055 ( .A(g11952), .ZN(g15055) );
INV_X32 U_g15065 ( .A(g12291), .ZN(g15065) );
INV_X32 U_g15074 ( .A(g11962), .ZN(g15074) );
INV_X32 U_g15080 ( .A(g12305), .ZN(g15080) );
INV_X32 U_I21415 ( .A(g11854), .ZN(I21415) );
INV_X32 U_g15092 ( .A(I21415), .ZN(g15092) );
INV_X32 U_I21420 ( .A(g13166), .ZN(I21420) );
INV_X32 U_g15095 ( .A(I21420), .ZN(g15095) );
INV_X32 U_g15096 ( .A(g11800), .ZN(g15096) );
INV_X32 U_I21426 ( .A(g11661), .ZN(I21426) );
INV_X32 U_g15106 ( .A(I21426), .ZN(g15106) );
INV_X32 U_I21429 ( .A(g13027), .ZN(I21429) );
INV_X32 U_g15109 ( .A(I21429), .ZN(g15109) );
INV_X32 U_I21432 ( .A(g13044), .ZN(I21432) );
INV_X32 U_g15112 ( .A(I21432), .ZN(g15112) );
INV_X32 U_I21435 ( .A(g11662), .ZN(I21435) );
INV_X32 U_g15115 ( .A(I21435), .ZN(g15115) );
INV_X32 U_g15118 ( .A(g11807), .ZN(g15118) );
INV_X32 U_g15128 ( .A(g12091), .ZN(g15128) );
INV_X32 U_g15129 ( .A(g12094), .ZN(g15129) );
INV_X32 U_I21443 ( .A(g12923), .ZN(I21443) );
INV_X32 U_g15130 ( .A(I21443), .ZN(g15130) );
INV_X32 U_I21446 ( .A(g13029), .ZN(I21446) );
INV_X32 U_g15133 ( .A(I21446), .ZN(g15133) );
INV_X32 U_I21449 ( .A(g13047), .ZN(I21449) );
INV_X32 U_g15136 ( .A(I21449), .ZN(g15136) );
INV_X32 U_I21452 ( .A(g13030), .ZN(I21452) );
INV_X32 U_g15139 ( .A(I21452), .ZN(g15139) );
INV_X32 U_g15144 ( .A(g12109), .ZN(g15144) );
INV_X32 U_I21458 ( .A(g13050), .ZN(I21458) );
INV_X32 U_g15145 ( .A(I21458), .ZN(g15145) );
INV_X32 U_I21461 ( .A(g13052), .ZN(I21461) );
INV_X32 U_g15148 ( .A(I21461), .ZN(g15148) );
INV_X32 U_g15151 ( .A(g12005), .ZN(g15151) );
INV_X32 U_g15161 ( .A(g12327), .ZN(g15161) );
INV_X32 U_g15170 ( .A(g12125), .ZN(g15170) );
INV_X32 U_g15174 ( .A(g12136), .ZN(g15174) );
INV_X32 U_g15175 ( .A(g12139), .ZN(g15175) );
INV_X32 U_g15176 ( .A(g12142), .ZN(g15176) );
INV_X32 U_g15177 ( .A(g12339), .ZN(g15177) );
INV_X32 U_I21476 ( .A(g11672), .ZN(I21476) );
INV_X32 U_g15179 ( .A(I21476), .ZN(g15179) );
INV_X32 U_I21479 ( .A(g13035), .ZN(I21479) );
INV_X32 U_g15182 ( .A(I21479), .ZN(g15182) );
INV_X32 U_I21482 ( .A(g13058), .ZN(I21482) );
INV_X32 U_g15185 ( .A(I21482), .ZN(g15185) );
INV_X32 U_g15188 ( .A(g11833), .ZN(g15188) );
INV_X32 U_I21488 ( .A(g11673), .ZN(I21488) );
INV_X32 U_g15198 ( .A(I21488), .ZN(g15198) );
INV_X32 U_I21491 ( .A(g13038), .ZN(I21491) );
INV_X32 U_g15201 ( .A(I21491), .ZN(g15201) );
INV_X32 U_I21494 ( .A(g13061), .ZN(I21494) );
INV_X32 U_g15204 ( .A(I21494), .ZN(g15204) );
INV_X32 U_I21497 ( .A(g11674), .ZN(I21497) );
INV_X32 U_g15207 ( .A(I21497), .ZN(g15207) );
INV_X32 U_g15210 ( .A(g11840), .ZN(g15210) );
INV_X32 U_g15220 ( .A(g12163), .ZN(g15220) );
INV_X32 U_g15221 ( .A(g12166), .ZN(g15221) );
INV_X32 U_I21505 ( .A(g12952), .ZN(I21505) );
INV_X32 U_g15222 ( .A(I21505), .ZN(g15222) );
INV_X32 U_I21508 ( .A(g13040), .ZN(I21508) );
INV_X32 U_g15225 ( .A(I21508), .ZN(g15225) );
INV_X32 U_I21511 ( .A(g13064), .ZN(I21511) );
INV_X32 U_g15228 ( .A(I21511), .ZN(g15228) );
INV_X32 U_I21514 ( .A(g13041), .ZN(I21514) );
INV_X32 U_g15231 ( .A(I21514), .ZN(g15231) );
INV_X32 U_g15236 ( .A(g12181), .ZN(g15236) );
INV_X32 U_I21520 ( .A(g13067), .ZN(I21520) );
INV_X32 U_g15237 ( .A(I21520), .ZN(g15237) );
INV_X32 U_I21523 ( .A(g13069), .ZN(I21523) );
INV_X32 U_g15240 ( .A(I21523), .ZN(g15240) );
INV_X32 U_I21531 ( .A(g11683), .ZN(I21531) );
INV_X32 U_g15248 ( .A(I21531), .ZN(g15248) );
INV_X32 U_I21534 ( .A(g13045), .ZN(I21534) );
INV_X32 U_g15251 ( .A(I21534), .ZN(g15251) );
INV_X32 U_I21537 ( .A(g13071), .ZN(I21537) );
INV_X32 U_g15254 ( .A(I21537), .ZN(g15254) );
INV_X32 U_g15260 ( .A(g12198), .ZN(g15260) );
INV_X32 U_g15261 ( .A(g12201), .ZN(g15261) );
INV_X32 U_g15262 ( .A(g12204), .ZN(g15262) );
INV_X32 U_g15263 ( .A(g12369), .ZN(g15263) );
INV_X32 U_I21548 ( .A(g11684), .ZN(I21548) );
INV_X32 U_g15265 ( .A(I21548), .ZN(g15265) );
INV_X32 U_I21551 ( .A(g13048), .ZN(I21551) );
INV_X32 U_g15268 ( .A(I21551), .ZN(g15268) );
INV_X32 U_I21554 ( .A(g13074), .ZN(I21554) );
INV_X32 U_g15271 ( .A(I21554), .ZN(g15271) );
INV_X32 U_g15274 ( .A(g11875), .ZN(g15274) );
INV_X32 U_I21560 ( .A(g11685), .ZN(I21560) );
INV_X32 U_g15284 ( .A(I21560), .ZN(g15284) );
INV_X32 U_I21563 ( .A(g13051), .ZN(I21563) );
INV_X32 U_g15287 ( .A(I21563), .ZN(g15287) );
INV_X32 U_I21566 ( .A(g13077), .ZN(I21566) );
INV_X32 U_g15290 ( .A(I21566), .ZN(g15290) );
INV_X32 U_I21569 ( .A(g11686), .ZN(I21569) );
INV_X32 U_g15293 ( .A(I21569), .ZN(g15293) );
INV_X32 U_g15296 ( .A(g11882), .ZN(g15296) );
INV_X32 U_g15306 ( .A(g12225), .ZN(g15306) );
INV_X32 U_g15307 ( .A(g12228), .ZN(g15307) );
INV_X32 U_I21577 ( .A(g12981), .ZN(I21577) );
INV_X32 U_g15308 ( .A(I21577), .ZN(g15308) );
INV_X32 U_I21580 ( .A(g13053), .ZN(I21580) );
INV_X32 U_g15311 ( .A(I21580), .ZN(g15311) );
INV_X32 U_I21583 ( .A(g13080), .ZN(I21583) );
INV_X32 U_g15314 ( .A(I21583), .ZN(g15314) );
INV_X32 U_I21586 ( .A(g13054), .ZN(I21586) );
INV_X32 U_g15317 ( .A(I21586), .ZN(g15317) );
INV_X32 U_g15322 ( .A(g12239), .ZN(g15322) );
INV_X32 U_g15323 ( .A(g12242), .ZN(g15323) );
INV_X32 U_I21595 ( .A(g11691), .ZN(I21595) );
INV_X32 U_g15326 ( .A(I21595), .ZN(g15326) );
INV_X32 U_I21598 ( .A(g13059), .ZN(I21598) );
INV_X32 U_g15329 ( .A(I21598), .ZN(g15329) );
INV_X32 U_I21601 ( .A(g13087), .ZN(I21601) );
INV_X32 U_g15332 ( .A(I21601), .ZN(g15332) );
INV_X32 U_I21609 ( .A(g11692), .ZN(I21609) );
INV_X32 U_g15340 ( .A(I21609), .ZN(g15340) );
INV_X32 U_I21612 ( .A(g13062), .ZN(I21612) );
INV_X32 U_g15343 ( .A(I21612), .ZN(g15343) );
INV_X32 U_I21615 ( .A(g13090), .ZN(I21615) );
INV_X32 U_g15346 ( .A(I21615), .ZN(g15346) );
INV_X32 U_g15352 ( .A(g12253), .ZN(g15352) );
INV_X32 U_g15353 ( .A(g12256), .ZN(g15353) );
INV_X32 U_g15354 ( .A(g12259), .ZN(g15354) );
INV_X32 U_g15355 ( .A(g12388), .ZN(g15355) );
INV_X32 U_I21626 ( .A(g11693), .ZN(I21626) );
INV_X32 U_g15357 ( .A(I21626), .ZN(g15357) );
INV_X32 U_I21629 ( .A(g13065), .ZN(I21629) );
INV_X32 U_g15360 ( .A(I21629), .ZN(g15360) );
INV_X32 U_I21632 ( .A(g13093), .ZN(I21632) );
INV_X32 U_g15363 ( .A(I21632), .ZN(g15363) );
INV_X32 U_g15366 ( .A(g11917), .ZN(g15366) );
INV_X32 U_I21638 ( .A(g11694), .ZN(I21638) );
INV_X32 U_g15376 ( .A(I21638), .ZN(g15376) );
INV_X32 U_I21641 ( .A(g13068), .ZN(I21641) );
INV_X32 U_g15379 ( .A(I21641), .ZN(g15379) );
INV_X32 U_I21644 ( .A(g13096), .ZN(I21644) );
INV_X32 U_g15382 ( .A(I21644), .ZN(g15382) );
INV_X32 U_I21647 ( .A(g11695), .ZN(I21647) );
INV_X32 U_g15385 ( .A(I21647), .ZN(g15385) );
INV_X32 U_g15390 ( .A(g12279), .ZN(g15390) );
INV_X32 U_I21655 ( .A(g11696), .ZN(I21655) );
INV_X32 U_g15393 ( .A(I21655), .ZN(g15393) );
INV_X32 U_I21658 ( .A(g13072), .ZN(I21658) );
INV_X32 U_g15396 ( .A(I21658), .ZN(g15396) );
INV_X32 U_I21661 ( .A(g13098), .ZN(I21661) );
INV_X32 U_g15399 ( .A(I21661), .ZN(g15399) );
INV_X32 U_I21666 ( .A(g13100), .ZN(I21666) );
INV_X32 U_g15404 ( .A(I21666), .ZN(g15404) );
INV_X32 U_g15408 ( .A(g12282), .ZN(g15408) );
INV_X32 U_g15409 ( .A(g12285), .ZN(g15409) );
INV_X32 U_I21674 ( .A(g11698), .ZN(I21674) );
INV_X32 U_g15412 ( .A(I21674), .ZN(g15412) );
INV_X32 U_I21677 ( .A(g13075), .ZN(I21677) );
INV_X32 U_g15415 ( .A(I21677), .ZN(g15415) );
INV_X32 U_I21680 ( .A(g13102), .ZN(I21680) );
INV_X32 U_g15418 ( .A(I21680), .ZN(g15418) );
INV_X32 U_I21688 ( .A(g11699), .ZN(I21688) );
INV_X32 U_g15426 ( .A(I21688), .ZN(g15426) );
INV_X32 U_I21691 ( .A(g13078), .ZN(I21691) );
INV_X32 U_g15429 ( .A(I21691), .ZN(g15429) );
INV_X32 U_I21694 ( .A(g13105), .ZN(I21694) );
INV_X32 U_g15432 ( .A(I21694), .ZN(g15432) );
INV_X32 U_g15438 ( .A(g12296), .ZN(g15438) );
INV_X32 U_g15439 ( .A(g12299), .ZN(g15439) );
INV_X32 U_g15440 ( .A(g12302), .ZN(g15440) );
INV_X32 U_g15441 ( .A(g12418), .ZN(g15441) );
INV_X32 U_I21705 ( .A(g11700), .ZN(I21705) );
INV_X32 U_g15443 ( .A(I21705), .ZN(g15443) );
INV_X32 U_I21708 ( .A(g13081), .ZN(I21708) );
INV_X32 U_g15446 ( .A(I21708), .ZN(g15446) );
INV_X32 U_I21711 ( .A(g13108), .ZN(I21711) );
INV_X32 U_g15449 ( .A(I21711), .ZN(g15449) );
INV_X32 U_g15458 ( .A(g12312), .ZN(g15458) );
INV_X32 U_I21720 ( .A(g11701), .ZN(I21720) );
INV_X32 U_g15461 ( .A(I21720), .ZN(g15461) );
INV_X32 U_I21723 ( .A(g13088), .ZN(I21723) );
INV_X32 U_g15464 ( .A(I21723), .ZN(g15464) );
INV_X32 U_I21726 ( .A(g13112), .ZN(I21726) );
INV_X32 U_g15467 ( .A(I21726), .ZN(g15467) );
INV_X32 U_I21730 ( .A(g13089), .ZN(I21730) );
INV_X32 U_g15471 ( .A(I21730), .ZN(g15471) );
INV_X32 U_g15474 ( .A(g12315), .ZN(g15474) );
INV_X32 U_I21736 ( .A(g11702), .ZN(I21736) );
INV_X32 U_g15477 ( .A(I21736), .ZN(g15477) );
INV_X32 U_I21739 ( .A(g13091), .ZN(I21739) );
INV_X32 U_g15480 ( .A(I21739), .ZN(g15480) );
INV_X32 U_I21742 ( .A(g13114), .ZN(I21742) );
INV_X32 U_g15483 ( .A(I21742), .ZN(g15483) );
INV_X32 U_I21747 ( .A(g13116), .ZN(I21747) );
INV_X32 U_g15488 ( .A(I21747), .ZN(g15488) );
INV_X32 U_g15492 ( .A(g12318), .ZN(g15492) );
INV_X32 U_g15493 ( .A(g12321), .ZN(g15493) );
INV_X32 U_I21755 ( .A(g11704), .ZN(I21755) );
INV_X32 U_g15496 ( .A(I21755), .ZN(g15496) );
INV_X32 U_I21758 ( .A(g13094), .ZN(I21758) );
INV_X32 U_g15499 ( .A(I21758), .ZN(g15499) );
INV_X32 U_I21761 ( .A(g13118), .ZN(I21761) );
INV_X32 U_g15502 ( .A(I21761), .ZN(g15502) );
INV_X32 U_I21769 ( .A(g11705), .ZN(I21769) );
INV_X32 U_g15510 ( .A(I21769), .ZN(g15510) );
INV_X32 U_I21772 ( .A(g13097), .ZN(I21772) );
INV_X32 U_g15513 ( .A(I21772), .ZN(g15513) );
INV_X32 U_I21775 ( .A(g13121), .ZN(I21775) );
INV_X32 U_g15516 ( .A(I21775), .ZN(g15516) );
INV_X32 U_I21780 ( .A(g13305), .ZN(I21780) );
INV_X32 U_g15521 ( .A(I21780), .ZN(g15521) );
INV_X32 U_g15524 ( .A(g12333), .ZN(g15524) );
INV_X32 U_g15525 ( .A(g12336), .ZN(g15525) );
INV_X32 U_I21787 ( .A(g11707), .ZN(I21787) );
INV_X32 U_g15528 ( .A(I21787), .ZN(g15528) );
INV_X32 U_I21790 ( .A(g13099), .ZN(I21790) );
INV_X32 U_g15531 ( .A(I21790), .ZN(g15531) );
INV_X32 U_I21793 ( .A(g13123), .ZN(I21793) );
INV_X32 U_g15534 ( .A(I21793), .ZN(g15534) );
INV_X32 U_I21796 ( .A(g11708), .ZN(I21796) );
INV_X32 U_g15537 ( .A(I21796), .ZN(g15537) );
INV_X32 U_g15544 ( .A(g12340), .ZN(g15544) );
INV_X32 U_I21803 ( .A(g11709), .ZN(I21803) );
INV_X32 U_g15547 ( .A(I21803), .ZN(g15547) );
INV_X32 U_I21806 ( .A(g13103), .ZN(I21806) );
INV_X32 U_g15550 ( .A(I21806), .ZN(g15550) );
INV_X32 U_I21809 ( .A(g13125), .ZN(I21809) );
INV_X32 U_g15553 ( .A(I21809), .ZN(g15553) );
INV_X32 U_I21813 ( .A(g13104), .ZN(I21813) );
INV_X32 U_g15557 ( .A(I21813), .ZN(g15557) );
INV_X32 U_g15560 ( .A(g12343), .ZN(g15560) );
INV_X32 U_I21819 ( .A(g11710), .ZN(I21819) );
INV_X32 U_g15563 ( .A(I21819), .ZN(g15563) );
INV_X32 U_I21822 ( .A(g13106), .ZN(I21822) );
INV_X32 U_g15566 ( .A(I21822), .ZN(g15566) );
INV_X32 U_I21825 ( .A(g13127), .ZN(I21825) );
INV_X32 U_g15569 ( .A(I21825), .ZN(g15569) );
INV_X32 U_I21830 ( .A(g13129), .ZN(I21830) );
INV_X32 U_g15574 ( .A(I21830), .ZN(g15574) );
INV_X32 U_g15578 ( .A(g12346), .ZN(g15578) );
INV_X32 U_g15579 ( .A(g12349), .ZN(g15579) );
INV_X32 U_I21838 ( .A(g11712), .ZN(I21838) );
INV_X32 U_g15582 ( .A(I21838), .ZN(g15582) );
INV_X32 U_I21841 ( .A(g13109), .ZN(I21841) );
INV_X32 U_g15585 ( .A(I21841), .ZN(g15585) );
INV_X32 U_I21844 ( .A(g13131), .ZN(I21844) );
INV_X32 U_g15588 ( .A(I21844), .ZN(g15588) );
INV_X32 U_I21852 ( .A(g11716), .ZN(I21852) );
INV_X32 U_g15596 ( .A(I21852), .ZN(g15596) );
INV_X32 U_I21855 ( .A(g13113), .ZN(I21855) );
INV_X32 U_g15599 ( .A(I21855), .ZN(g15599) );
INV_X32 U_g15602 ( .A(g12363), .ZN(g15602) );
INV_X32 U_g15603 ( .A(g12366), .ZN(g15603) );
INV_X32 U_I21862 ( .A(g11717), .ZN(I21862) );
INV_X32 U_g15606 ( .A(I21862), .ZN(g15606) );
INV_X32 U_I21865 ( .A(g13115), .ZN(I21865) );
INV_X32 U_g15609 ( .A(I21865), .ZN(g15609) );
INV_X32 U_I21868 ( .A(g13134), .ZN(I21868) );
INV_X32 U_g15612 ( .A(I21868), .ZN(g15612) );
INV_X32 U_I21871 ( .A(g11718), .ZN(I21871) );
INV_X32 U_g15615 ( .A(I21871), .ZN(g15615) );
INV_X32 U_g15622 ( .A(g12370), .ZN(g15622) );
INV_X32 U_I21878 ( .A(g11719), .ZN(I21878) );
INV_X32 U_g15625 ( .A(I21878), .ZN(g15625) );
INV_X32 U_I21881 ( .A(g13119), .ZN(I21881) );
INV_X32 U_g15628 ( .A(I21881), .ZN(g15628) );
INV_X32 U_I21884 ( .A(g13136), .ZN(I21884) );
INV_X32 U_g15631 ( .A(I21884), .ZN(g15631) );
INV_X32 U_I21888 ( .A(g13120), .ZN(I21888) );
INV_X32 U_g15635 ( .A(I21888), .ZN(g15635) );
INV_X32 U_g15638 ( .A(g12373), .ZN(g15638) );
INV_X32 U_I21894 ( .A(g11720), .ZN(I21894) );
INV_X32 U_g15641 ( .A(I21894), .ZN(g15641) );
INV_X32 U_I21897 ( .A(g13122), .ZN(I21897) );
INV_X32 U_g15644 ( .A(I21897), .ZN(g15644) );
INV_X32 U_I21900 ( .A(g13138), .ZN(I21900) );
INV_X32 U_g15647 ( .A(I21900), .ZN(g15647) );
INV_X32 U_I21905 ( .A(g13140), .ZN(I21905) );
INV_X32 U_g15652 ( .A(I21905), .ZN(g15652) );
INV_X32 U_I21908 ( .A(g13082), .ZN(I21908) );
INV_X32 U_g15655 ( .A(I21908), .ZN(g15655) );
INV_X32 U_g15659 ( .A(g11706), .ZN(g15659) );
INV_X32 U_g15665 ( .A(g12379), .ZN(g15665) );
INV_X32 U_I21918 ( .A(g11721), .ZN(I21918) );
INV_X32 U_g15667 ( .A(I21918), .ZN(g15667) );
INV_X32 U_I21923 ( .A(g11722), .ZN(I21923) );
INV_X32 U_g15672 ( .A(I21923), .ZN(g15672) );
INV_X32 U_I21926 ( .A(g13126), .ZN(I21926) );
INV_X32 U_g15675 ( .A(I21926), .ZN(g15675) );
INV_X32 U_g15678 ( .A(g12382), .ZN(g15678) );
INV_X32 U_g15679 ( .A(g12385), .ZN(g15679) );
INV_X32 U_I21933 ( .A(g11723), .ZN(I21933) );
INV_X32 U_g15682 ( .A(I21933), .ZN(g15682) );
INV_X32 U_I21936 ( .A(g13128), .ZN(I21936) );
INV_X32 U_g15685 ( .A(I21936), .ZN(g15685) );
INV_X32 U_I21939 ( .A(g13142), .ZN(I21939) );
INV_X32 U_g15688 ( .A(I21939), .ZN(g15688) );
INV_X32 U_I21942 ( .A(g11724), .ZN(I21942) );
INV_X32 U_g15691 ( .A(I21942), .ZN(g15691) );
INV_X32 U_g15698 ( .A(g12389), .ZN(g15698) );
INV_X32 U_I21949 ( .A(g11725), .ZN(I21949) );
INV_X32 U_g15701 ( .A(I21949), .ZN(g15701) );
INV_X32 U_I21952 ( .A(g13132), .ZN(I21952) );
INV_X32 U_g15704 ( .A(I21952), .ZN(g15704) );
INV_X32 U_I21955 ( .A(g13144), .ZN(I21955) );
INV_X32 U_g15707 ( .A(I21955), .ZN(g15707) );
INV_X32 U_I21959 ( .A(g13133), .ZN(I21959) );
INV_X32 U_g15711 ( .A(I21959), .ZN(g15711) );
INV_X32 U_I21962 ( .A(g13004), .ZN(I21962) );
INV_X32 U_g15714 ( .A(I21962), .ZN(g15714) );
INV_X32 U_g15722 ( .A(g13011), .ZN(g15722) );
INV_X32 U_g15724 ( .A(g12409), .ZN(g15724) );
INV_X32 U_I21974 ( .A(g11726), .ZN(I21974) );
INV_X32 U_g15726 ( .A(I21974), .ZN(g15726) );
INV_X32 U_I21979 ( .A(g11727), .ZN(I21979) );
INV_X32 U_g15731 ( .A(I21979), .ZN(g15731) );
INV_X32 U_I21982 ( .A(g13137), .ZN(I21982) );
INV_X32 U_g15734 ( .A(I21982), .ZN(g15734) );
INV_X32 U_g15737 ( .A(g12412), .ZN(g15737) );
INV_X32 U_g15738 ( .A(g12415), .ZN(g15738) );
INV_X32 U_I21989 ( .A(g11728), .ZN(I21989) );
INV_X32 U_g15741 ( .A(I21989), .ZN(g15741) );
INV_X32 U_I21992 ( .A(g13139), .ZN(I21992) );
INV_X32 U_g15744 ( .A(I21992), .ZN(g15744) );
INV_X32 U_I21995 ( .A(g13146), .ZN(I21995) );
INV_X32 U_g15747 ( .A(I21995), .ZN(g15747) );
INV_X32 U_I21998 ( .A(g11729), .ZN(I21998) );
INV_X32 U_g15750 ( .A(I21998), .ZN(g15750) );
INV_X32 U_g15762 ( .A(g13011), .ZN(g15762) );
INV_X32 U_g15764 ( .A(g12421), .ZN(g15764) );
INV_X32 U_I22014 ( .A(g11730), .ZN(I22014) );
INV_X32 U_g15766 ( .A(I22014), .ZN(g15766) );
INV_X32 U_I22019 ( .A(g11731), .ZN(I22019) );
INV_X32 U_g15771 ( .A(I22019), .ZN(g15771) );
INV_X32 U_I22022 ( .A(g13145), .ZN(I22022) );
INV_X32 U_g15774 ( .A(I22022), .ZN(g15774) );
INV_X32 U_I22025 ( .A(g11617), .ZN(I22025) );
INV_X32 U_g15777 ( .A(I22025), .ZN(g15777) );
INV_X32 U_g15790 ( .A(g13011), .ZN(g15790) );
INV_X32 U_g15792 ( .A(g12426), .ZN(g15792) );
INV_X32 U_I22044 ( .A(g11733), .ZN(I22044) );
INV_X32 U_g15794 ( .A(I22044), .ZN(g15794) );
INV_X32 U_g15800 ( .A(g12909), .ZN(g15800) );
INV_X32 U_g15813 ( .A(g13011), .ZN(g15813) );
INV_X32 U_g15859 ( .A(g13378), .ZN(g15859) );
INV_X32 U_I22120 ( .A(g12909), .ZN(I22120) );
INV_X32 U_g15876 ( .A(I22120), .ZN(g15876) );
INV_X32 U_g15880 ( .A(g11624), .ZN(g15880) );
INV_X32 U_g15890 ( .A(g11600), .ZN(g15890) );
INV_X32 U_g15904 ( .A(g11644), .ZN(g15904) );
INV_X32 U_g15913 ( .A(g11647), .ZN(g15913) );
INV_X32 U_g15923 ( .A(g11630), .ZN(g15923) );
INV_X32 U_g15933 ( .A(g11663), .ZN(g15933) );
INV_X32 U_g15942 ( .A(g11666), .ZN(g15942) );
INV_X32 U_g15952 ( .A(g11653), .ZN(g15952) );
INV_X32 U_g15962 ( .A(g11675), .ZN(g15962) );
INV_X32 U_g15971 ( .A(g11678), .ZN(g15971) );
INV_X32 U_g15981 ( .A(g11687), .ZN(g15981) );
INV_X32 U_I22163 ( .A(g12433), .ZN(I22163) );
INV_X32 U_g15989 ( .A(I22163), .ZN(g15989) );
INV_X32 U_g15991 ( .A(g12548), .ZN(g15991) );
INV_X32 U_g15994 ( .A(g12555), .ZN(g15994) );
INV_X32 U_g15997 ( .A(g12561), .ZN(g15997) );
INV_X32 U_g16001 ( .A(g12601), .ZN(g16001) );
INV_X32 U_g16002 ( .A(g12604), .ZN(g16002) );
INV_X32 U_g16005 ( .A(g12608), .ZN(g16005) );
INV_X32 U_g16007 ( .A(g12647), .ZN(g16007) );
INV_X32 U_g16011 ( .A(g12651), .ZN(g16011) );
INV_X32 U_g16012 ( .A(g12654), .ZN(g16012) );
INV_X32 U_g16013 ( .A(g12692), .ZN(g16013) );
INV_X32 U_g16014 ( .A(g12695), .ZN(g16014) );
INV_X32 U_g16023 ( .A(g12699), .ZN(g16023) );
INV_X32 U_g16024 ( .A(g12702), .ZN(g16024) );
INV_X32 U_g16025 ( .A(g12705), .ZN(g16025) );
INV_X32 U_g16026 ( .A(g12708), .ZN(g16026) );
INV_X32 U_g16027 ( .A(g12744), .ZN(g16027) );
INV_X32 U_g16034 ( .A(g12749), .ZN(g16034) );
INV_X32 U_g16035 ( .A(g12752), .ZN(g16035) );
INV_X32 U_g16039 ( .A(g12756), .ZN(g16039) );
INV_X32 U_g16040 ( .A(g12759), .ZN(g16040) );
INV_X32 U_g16041 ( .A(g12762), .ZN(g16041) );
INV_X32 U_g16042 ( .A(g12765), .ZN(g16042) );
INV_X32 U_g16043 ( .A(g12769), .ZN(g16043) );
INV_X32 U_g16044 ( .A(g12772), .ZN(g16044) );
INV_X32 U_g16054 ( .A(g12783), .ZN(g16054) );
INV_X32 U_g16055 ( .A(g12786), .ZN(g16055) );
INV_X32 U_g16056 ( .A(g12791), .ZN(g16056) );
INV_X32 U_g16057 ( .A(g12794), .ZN(g16057) );
INV_X32 U_g16061 ( .A(g12798), .ZN(g16061) );
INV_X32 U_g16062 ( .A(g12801), .ZN(g16062) );
INV_X32 U_g16063 ( .A(g12804), .ZN(g16063) );
INV_X32 U_g16064 ( .A(g12808), .ZN(g16064) );
INV_X32 U_g16065 ( .A(g12811), .ZN(g16065) );
INV_X32 U_g16075 ( .A(g11861), .ZN(g16075) );
INV_X32 U_g16088 ( .A(g12816), .ZN(g16088) );
INV_X32 U_g16090 ( .A(g12822), .ZN(g16090) );
INV_X32 U_g16091 ( .A(g12825), .ZN(g16091) );
INV_X32 U_g16092 ( .A(g12830), .ZN(g16092) );
INV_X32 U_g16093 ( .A(g12833), .ZN(g16093) );
INV_X32 U_g16097 ( .A(g12837), .ZN(g16097) );
INV_X32 U_g16098 ( .A(g12840), .ZN(g16098) );
INV_X32 U_g16099 ( .A(g12844), .ZN(g16099) );
INV_X32 U_g16113 ( .A(g11903), .ZN(g16113) );
INV_X32 U_g16126 ( .A(g12854), .ZN(g16126) );
INV_X32 U_g16128 ( .A(g12860), .ZN(g16128) );
INV_X32 U_g16129 ( .A(g12863), .ZN(g16129) );
INV_X32 U_g16130 ( .A(g12868), .ZN(g16130) );
INV_X32 U_g16131 ( .A(g12871), .ZN(g16131) );
INV_X32 U_g16142 ( .A(g13057), .ZN(g16142) );
INV_X32 U_g16154 ( .A(g12194), .ZN(g16154) );
INV_X32 U_g16164 ( .A(g11953), .ZN(g16164) );
INV_X32 U_g16177 ( .A(g12895), .ZN(g16177) );
INV_X32 U_g16179 ( .A(g12901), .ZN(g16179) );
INV_X32 U_g16180 ( .A(g12904), .ZN(g16180) );
INV_X32 U_g16189 ( .A(g13043), .ZN(g16189) );
INV_X32 U_g16201 ( .A(g13073), .ZN(g16201) );
INV_X32 U_g16213 ( .A(g12249), .ZN(g16213) );
INV_X32 U_g16223 ( .A(g12006), .ZN(g16223) );
INV_X32 U_g16236 ( .A(g12935), .ZN(g16236) );
INV_X32 U_g16243 ( .A(g13033), .ZN(g16243) );
INV_X32 U_g16254 ( .A(g13060), .ZN(g16254) );
INV_X32 U_g16266 ( .A(g13092), .ZN(g16266) );
INV_X32 U_g16278 ( .A(g12292), .ZN(g16278) );
INV_X32 U_g16287 ( .A(g12962), .ZN(g16287) );
INV_X32 U_g16293 ( .A(g13025), .ZN(g16293) );
INV_X32 U_I22382 ( .A(g520), .ZN(I22382) );
INV_X32 U_g16297 ( .A(I22382), .ZN(g16297) );
INV_X32 U_g16302 ( .A(g13046), .ZN(g16302) );
INV_X32 U_g16313 ( .A(g13076), .ZN(g16313) );
INV_X32 U_g16325 ( .A(g13107), .ZN(g16325) );
INV_X32 U_g16337 ( .A(g12328), .ZN(g16337) );
INV_X32 U_g16351 ( .A(g13036), .ZN(g16351) );
INV_X32 U_I22414 ( .A(g1206), .ZN(I22414) );
INV_X32 U_g16355 ( .A(I22414), .ZN(g16355) );
INV_X32 U_g16360 ( .A(g13063), .ZN(g16360) );
INV_X32 U_g16371 ( .A(g13095), .ZN(g16371) );
INV_X32 U_g16395 ( .A(g13049), .ZN(g16395) );
INV_X32 U_I22444 ( .A(g1900), .ZN(I22444) );
INV_X32 U_g16399 ( .A(I22444), .ZN(g16399) );
INV_X32 U_g16404 ( .A(g13079), .ZN(g16404) );
INV_X32 U_g16433 ( .A(g13066), .ZN(g16433) );
INV_X32 U_I22475 ( .A(g2594), .ZN(I22475) );
INV_X32 U_g16437 ( .A(I22475), .ZN(g16437) );
INV_X32 U_g16466 ( .A(g12017), .ZN(g16466) );
INV_X32 U_I22503 ( .A(g13598), .ZN(I22503) );
INV_X32 U_g16467 ( .A(I22503), .ZN(g16467) );
INV_X32 U_I22506 ( .A(g13624), .ZN(I22506) );
INV_X32 U_g16468 ( .A(I22506), .ZN(g16468) );
INV_X32 U_I22509 ( .A(g13610), .ZN(I22509) );
INV_X32 U_g16469 ( .A(I22509), .ZN(g16469) );
INV_X32 U_I22512 ( .A(g13635), .ZN(I22512) );
INV_X32 U_g16470 ( .A(I22512), .ZN(g16470) );
INV_X32 U_I22515 ( .A(g13620), .ZN(I22515) );
INV_X32 U_g16471 ( .A(I22515), .ZN(g16471) );
INV_X32 U_I22518 ( .A(g13647), .ZN(I22518) );
INV_X32 U_g16472 ( .A(I22518), .ZN(g16472) );
INV_X32 U_I22521 ( .A(g13632), .ZN(I22521) );
INV_X32 U_g16473 ( .A(I22521), .ZN(g16473) );
INV_X32 U_I22524 ( .A(g13673), .ZN(I22524) );
INV_X32 U_g16474 ( .A(I22524), .ZN(g16474) );
INV_X32 U_I22527 ( .A(g13469), .ZN(I22527) );
INV_X32 U_g16475 ( .A(I22527), .ZN(g16475) );
INV_X32 U_I22530 ( .A(g14774), .ZN(I22530) );
INV_X32 U_g16476 ( .A(I22530), .ZN(g16476) );
INV_X32 U_I22533 ( .A(g14795), .ZN(I22533) );
INV_X32 U_g16477 ( .A(I22533), .ZN(g16477) );
INV_X32 U_I22536 ( .A(g14829), .ZN(I22536) );
INV_X32 U_g16478 ( .A(I22536), .ZN(g16478) );
INV_X32 U_I22539 ( .A(g14882), .ZN(I22539) );
INV_X32 U_g16479 ( .A(I22539), .ZN(g16479) );
INV_X32 U_I22542 ( .A(g14954), .ZN(I22542) );
INV_X32 U_g16480 ( .A(I22542), .ZN(g16480) );
INV_X32 U_I22545 ( .A(g15018), .ZN(I22545) );
INV_X32 U_g16481 ( .A(I22545), .ZN(g16481) );
INV_X32 U_I22548 ( .A(g14718), .ZN(I22548) );
INV_X32 U_g16482 ( .A(I22548), .ZN(g16482) );
INV_X32 U_I22551 ( .A(g14745), .ZN(I22551) );
INV_X32 U_g16483 ( .A(I22551), .ZN(g16483) );
INV_X32 U_I22554 ( .A(g14765), .ZN(I22554) );
INV_X32 U_g16484 ( .A(I22554), .ZN(g16484) );
INV_X32 U_I22557 ( .A(g14775), .ZN(I22557) );
INV_X32 U_g16485 ( .A(I22557), .ZN(g16485) );
INV_X32 U_I22560 ( .A(g14796), .ZN(I22560) );
INV_X32 U_g16486 ( .A(I22560), .ZN(g16486) );
INV_X32 U_I22563 ( .A(g14830), .ZN(I22563) );
INV_X32 U_g16487 ( .A(I22563), .ZN(g16487) );
INV_X32 U_I22566 ( .A(g14883), .ZN(I22566) );
INV_X32 U_g16488 ( .A(I22566), .ZN(g16488) );
INV_X32 U_I22569 ( .A(g14955), .ZN(I22569) );
INV_X32 U_g16489 ( .A(I22569), .ZN(g16489) );
INV_X32 U_I22572 ( .A(g15019), .ZN(I22572) );
INV_X32 U_g16490 ( .A(I22572), .ZN(g16490) );
INV_X32 U_I22575 ( .A(g15092), .ZN(I22575) );
INV_X32 U_g16491 ( .A(I22575), .ZN(g16491) );
INV_X32 U_I22578 ( .A(g14746), .ZN(I22578) );
INV_X32 U_g16492 ( .A(I22578), .ZN(g16492) );
INV_X32 U_I22581 ( .A(g14766), .ZN(I22581) );
INV_X32 U_g16493 ( .A(I22581), .ZN(g16493) );
INV_X32 U_I22584 ( .A(g15989), .ZN(I22584) );
INV_X32 U_g16494 ( .A(I22584), .ZN(g16494) );
INV_X32 U_I22587 ( .A(g14684), .ZN(I22587) );
INV_X32 U_g16495 ( .A(I22587), .ZN(g16495) );
INV_X32 U_I22590 ( .A(g13863), .ZN(I22590) );
INV_X32 U_g16496 ( .A(I22590), .ZN(g16496) );
INV_X32 U_I22593 ( .A(g15876), .ZN(I22593) );
INV_X32 U_g16497 ( .A(I22593), .ZN(g16497) );
INV_X32 U_g16501 ( .A(g14158), .ZN(g16501) );
INV_X32 U_I22599 ( .A(g14966), .ZN(I22599) );
INV_X32 U_g16506 ( .A(I22599), .ZN(g16506) );
INV_X32 U_g16507 ( .A(g14186), .ZN(g16507) );
INV_X32 U_I22604 ( .A(g15080), .ZN(I22604) );
INV_X32 U_g16514 ( .A(I22604), .ZN(g16514) );
INV_X32 U_g16515 ( .A(g14244), .ZN(g16515) );
INV_X32 U_g16523 ( .A(g14273), .ZN(g16523) );
INV_X32 U_I22611 ( .A(g15055), .ZN(I22611) );
INV_X32 U_g16528 ( .A(I22611), .ZN(g16528) );
INV_X32 U_g16529 ( .A(g14301), .ZN(g16529) );
INV_X32 U_I22618 ( .A(g14630), .ZN(I22618) );
INV_X32 U_g16540 ( .A(I22618), .ZN(g16540) );
INV_X32 U_g16543 ( .A(g14347), .ZN(g16543) );
INV_X32 U_g16546 ( .A(g14366), .ZN(g16546) );
INV_X32 U_g16554 ( .A(g14395), .ZN(g16554) );
INV_X32 U_I22626 ( .A(g15151), .ZN(I22626) );
INV_X32 U_g16559 ( .A(I22626), .ZN(g16559) );
INV_X32 U_g16560 ( .A(g14423), .ZN(g16560) );
INV_X32 U_I22640 ( .A(g14650), .ZN(I22640) );
INV_X32 U_g16572 ( .A(I22640), .ZN(g16572) );
INV_X32 U_g16575 ( .A(g14459), .ZN(g16575) );
INV_X32 U_g16578 ( .A(g14478), .ZN(g16578) );
INV_X32 U_g16586 ( .A(g14507), .ZN(g16586) );
INV_X32 U_I22651 ( .A(g14677), .ZN(I22651) );
INV_X32 U_g16596 ( .A(I22651), .ZN(g16596) );
INV_X32 U_g16599 ( .A(g14546), .ZN(g16599) );
INV_X32 U_g16602 ( .A(g14565), .ZN(g16602) );
INV_X32 U_I22657 ( .A(g14657), .ZN(I22657) );
INV_X32 U_g16608 ( .A(I22657), .ZN(g16608) );
INV_X32 U_I22663 ( .A(g14711), .ZN(I22663) );
INV_X32 U_g16616 ( .A(I22663), .ZN(g16616) );
INV_X32 U_g16619 ( .A(g14601), .ZN(g16619) );
INV_X32 U_I22667 ( .A(g14642), .ZN(I22667) );
INV_X32 U_g16622 ( .A(I22667), .ZN(g16622) );
INV_X32 U_I22671 ( .A(g14691), .ZN(I22671) );
INV_X32 U_g16626 ( .A(I22671), .ZN(g16626) );
INV_X32 U_I22676 ( .A(g14630), .ZN(I22676) );
INV_X32 U_g16633 ( .A(I22676), .ZN(g16633) );
INV_X32 U_I22679 ( .A(g14669), .ZN(I22679) );
INV_X32 U_g16636 ( .A(I22679), .ZN(g16636) );
INV_X32 U_I22683 ( .A(g14725), .ZN(I22683) );
INV_X32 U_g16640 ( .A(I22683), .ZN(g16640) );
INV_X32 U_I22687 ( .A(g14650), .ZN(I22687) );
INV_X32 U_g16644 ( .A(I22687), .ZN(g16644) );
INV_X32 U_I22690 ( .A(g14703), .ZN(I22690) );
INV_X32 U_g16647 ( .A(I22690), .ZN(g16647) );
INV_X32 U_I22694 ( .A(g14753), .ZN(I22694) );
INV_X32 U_g16651 ( .A(I22694), .ZN(g16651) );
INV_X32 U_I22699 ( .A(g14677), .ZN(I22699) );
INV_X32 U_g16656 ( .A(I22699), .ZN(g16656) );
INV_X32 U_I22702 ( .A(g14737), .ZN(I22702) );
INV_X32 U_g16659 ( .A(I22702), .ZN(g16659) );
INV_X32 U_g16665 ( .A(g14776), .ZN(g16665) );
INV_X32 U_I22715 ( .A(g14711), .ZN(I22715) );
INV_X32 U_g16673 ( .A(I22715), .ZN(g16673) );
INV_X32 U_I22718 ( .A(g14657), .ZN(I22718) );
INV_X32 U_g16676 ( .A(I22718), .ZN(g16676) );
INV_X32 U_g16682 ( .A(g14797), .ZN(g16682) );
INV_X32 U_g16686 ( .A(g14811), .ZN(g16686) );
INV_X32 U_I22726 ( .A(g14642), .ZN(I22726) );
INV_X32 U_g16694 ( .A(I22726), .ZN(g16694) );
INV_X32 U_g16697 ( .A(g14837), .ZN(g16697) );
INV_X32 U_I22730 ( .A(g14691), .ZN(I22730) );
INV_X32 U_g16702 ( .A(I22730), .ZN(g16702) );
INV_X32 U_g16708 ( .A(g14849), .ZN(g16708) );
INV_X32 U_g16712 ( .A(g14863), .ZN(g16712) );
INV_X32 U_I22737 ( .A(g14630), .ZN(I22737) );
INV_X32 U_g16719 ( .A(I22737), .ZN(g16719) );
INV_X32 U_g16722 ( .A(g14895), .ZN(g16722) );
INV_X32 U_I22741 ( .A(g14669), .ZN(I22741) );
INV_X32 U_g16725 ( .A(I22741), .ZN(g16725) );
INV_X32 U_g16728 ( .A(g14910), .ZN(g16728) );
INV_X32 U_I22745 ( .A(g14725), .ZN(I22745) );
INV_X32 U_g16733 ( .A(I22745), .ZN(g16733) );
INV_X32 U_g16739 ( .A(g14922), .ZN(g16739) );
INV_X32 U_g16743 ( .A(g14936), .ZN(g16743) );
INV_X32 U_g16749 ( .A(g15782), .ZN(g16749) );
INV_X32 U_I22752 ( .A(g14657), .ZN(I22752) );
INV_X32 U_g16758 ( .A(I22752), .ZN(g16758) );
INV_X32 U_I22755 ( .A(g14650), .ZN(I22755) );
INV_X32 U_g16761 ( .A(I22755), .ZN(g16761) );
INV_X32 U_g16764 ( .A(g14976), .ZN(g16764) );
INV_X32 U_I22759 ( .A(g14703), .ZN(I22759) );
INV_X32 U_g16767 ( .A(I22759), .ZN(g16767) );
INV_X32 U_g16770 ( .A(g14991), .ZN(g16770) );
INV_X32 U_I22763 ( .A(g14753), .ZN(I22763) );
INV_X32 U_g16775 ( .A(I22763), .ZN(g16775) );
INV_X32 U_g16781 ( .A(g15003), .ZN(g16781) );
INV_X32 U_I22768 ( .A(g14691), .ZN(I22768) );
INV_X32 U_g16785 ( .A(I22768), .ZN(g16785) );
INV_X32 U_I22771 ( .A(g14677), .ZN(I22771) );
INV_X32 U_g16788 ( .A(I22771), .ZN(g16788) );
INV_X32 U_g16791 ( .A(g15065), .ZN(g16791) );
INV_X32 U_I22775 ( .A(g14737), .ZN(I22775) );
INV_X32 U_g16794 ( .A(I22775), .ZN(g16794) );
INV_X32 U_g16797 ( .A(g15080), .ZN(g16797) );
INV_X32 U_g16804 ( .A(g15803), .ZN(g16804) );
INV_X32 U_g16809 ( .A(g15842), .ZN(g16809) );
INV_X32 U_I22783 ( .A(g13572), .ZN(I22783) );
INV_X32 U_g16813 ( .A(I22783), .ZN(g16813) );
INV_X32 U_I22786 ( .A(g14725), .ZN(I22786) );
INV_X32 U_g16814 ( .A(I22786), .ZN(g16814) );
INV_X32 U_I22789 ( .A(g14711), .ZN(I22789) );
INV_X32 U_g16817 ( .A(I22789), .ZN(g16817) );
INV_X32 U_g16820 ( .A(g15161), .ZN(g16820) );
INV_X32 U_g16825 ( .A(g15855), .ZN(g16825) );
INV_X32 U_I22797 ( .A(g14165), .ZN(I22797) );
INV_X32 U_g16830 ( .A(I22797), .ZN(g16830) );
INV_X32 U_I22800 ( .A(g13581), .ZN(I22800) );
INV_X32 U_g16831 ( .A(I22800), .ZN(g16831) );
INV_X32 U_I22803 ( .A(g14753), .ZN(I22803) );
INV_X32 U_g16832 ( .A(I22803), .ZN(g16832) );
INV_X32 U_g16836 ( .A(g15818), .ZN(g16836) );
INV_X32 U_g16840 ( .A(g15878), .ZN(g16840) );
INV_X32 U_I22810 ( .A(g14280), .ZN(I22810) );
INV_X32 U_g16842 ( .A(I22810), .ZN(g16842) );
INV_X32 U_I22813 ( .A(g13601), .ZN(I22813) );
INV_X32 U_g16843 ( .A(I22813), .ZN(g16843) );
INV_X32 U_g16846 ( .A(g15903), .ZN(g16846) );
INV_X32 U_I22820 ( .A(g14402), .ZN(I22820) );
INV_X32 U_g16848 ( .A(I22820), .ZN(g16848) );
INV_X32 U_I22823 ( .A(g13613), .ZN(I22823) );
INV_X32 U_g16849 ( .A(I22823), .ZN(g16849) );
INV_X32 U_I22828 ( .A(g14514), .ZN(I22828) );
INV_X32 U_g16852 ( .A(I22828), .ZN(g16852) );
INV_X32 U_I22836 ( .A(g13571), .ZN(I22836) );
INV_X32 U_g16858 ( .A(I22836), .ZN(g16858) );
INV_X32 U_I22842 ( .A(g13580), .ZN(I22842) );
INV_X32 U_g16862 ( .A(I22842), .ZN(g16862) );
INV_X32 U_I22845 ( .A(g13579), .ZN(I22845) );
INV_X32 U_g16863 ( .A(I22845), .ZN(g16863) );
INV_X32 U_g16867 ( .A(g13589), .ZN(g16867) );
INV_X32 U_I22852 ( .A(g13600), .ZN(I22852) );
INV_X32 U_g16877 ( .A(I22852), .ZN(g16877) );
INV_X32 U_I22855 ( .A(g13588), .ZN(I22855) );
INV_X32 U_g16878 ( .A(I22855), .ZN(g16878) );
INV_X32 U_I22860 ( .A(g14885), .ZN(I22860) );
INV_X32 U_g16881 ( .A(I22860), .ZN(g16881) );
INV_X32 U_g16884 ( .A(g13589), .ZN(g16884) );
INV_X32 U_g16895 ( .A(g13589), .ZN(g16895) );
INV_X32 U_I22866 ( .A(g13612), .ZN(I22866) );
INV_X32 U_g16905 ( .A(I22866), .ZN(g16905) );
INV_X32 U_I22869 ( .A(g13608), .ZN(I22869) );
INV_X32 U_g16906 ( .A(I22869), .ZN(g16906) );
INV_X32 U_I22875 ( .A(g14966), .ZN(I22875) );
INV_X32 U_g16910 ( .A(I22875), .ZN(g16910) );
INV_X32 U_g16913 ( .A(g13589), .ZN(g16913) );
INV_X32 U_g16924 ( .A(g13589), .ZN(g16924) );
INV_X32 U_I22881 ( .A(g13622), .ZN(I22881) );
INV_X32 U_g16934 ( .A(I22881), .ZN(g16934) );
INV_X32 U_I22893 ( .A(g15055), .ZN(I22893) );
INV_X32 U_g16940 ( .A(I22893), .ZN(g16940) );
INV_X32 U_g16943 ( .A(g13589), .ZN(g16943) );
INV_X32 U_g16954 ( .A(g13589), .ZN(g16954) );
INV_X32 U_I22912 ( .A(g15151), .ZN(I22912) );
INV_X32 U_g16971 ( .A(I22912), .ZN(g16971) );
INV_X32 U_g16974 ( .A(g13589), .ZN(g16974) );
INV_X32 U_g17029 ( .A(g14685), .ZN(g17029) );
INV_X32 U_g17057 ( .A(g13519), .ZN(g17057) );
INV_X32 U_g17063 ( .A(g14719), .ZN(g17063) );
INV_X32 U_g17092 ( .A(g13530), .ZN(g17092) );
INV_X32 U_g17098 ( .A(g14747), .ZN(g17098) );
INV_X32 U_g17130 ( .A(g13541), .ZN(g17130) );
INV_X32 U_g17136 ( .A(g14768), .ZN(g17136) );
INV_X32 U_g17157 ( .A(g13552), .ZN(g17157) );
INV_X32 U_I23253 ( .A(g13741), .ZN(I23253) );
INV_X32 U_g17189 ( .A(I23253), .ZN(g17189) );
INV_X32 U_I23274 ( .A(g13741), .ZN(I23274) );
INV_X32 U_g17200 ( .A(I23274), .ZN(g17200) );
INV_X32 U_g17203 ( .A(g13568), .ZN(g17203) );
INV_X32 U_I23287 ( .A(g13741), .ZN(I23287) );
INV_X32 U_g17207 ( .A(I23287), .ZN(g17207) );
INV_X32 U_g17208 ( .A(g13576), .ZN(g17208) );
INV_X32 U_I23292 ( .A(g13741), .ZN(I23292) );
INV_X32 U_g17212 ( .A(I23292), .ZN(g17212) );
INV_X32 U_g17214 ( .A(g13585), .ZN(g17214) );
INV_X32 U_g17217 ( .A(g13605), .ZN(g17217) );
INV_X32 U_I23309 ( .A(g16132), .ZN(I23309) );
INV_X32 U_g17227 ( .A(I23309), .ZN(g17227) );
INV_X32 U_I23314 ( .A(g15720), .ZN(I23314) );
INV_X32 U_g17230 ( .A(I23314), .ZN(g17230) );
INV_X32 U_I23317 ( .A(g16181), .ZN(I23317) );
INV_X32 U_g17233 ( .A(I23317), .ZN(g17233) );
INV_X32 U_I23323 ( .A(g15664), .ZN(I23323) );
INV_X32 U_g17237 ( .A(I23323), .ZN(g17237) );
INV_X32 U_I23326 ( .A(g15758), .ZN(I23326) );
INV_X32 U_g17240 ( .A(I23326), .ZN(g17240) );
INV_X32 U_I23329 ( .A(g15760), .ZN(I23329) );
INV_X32 U_g17243 ( .A(I23329), .ZN(g17243) );
INV_X32 U_I23335 ( .A(g16412), .ZN(I23335) );
INV_X32 U_g17249 ( .A(I23335), .ZN(g17249) );
INV_X32 U_I23338 ( .A(g15721), .ZN(I23338) );
INV_X32 U_g17252 ( .A(I23338), .ZN(g17252) );
INV_X32 U_I23341 ( .A(g15784), .ZN(I23341) );
INV_X32 U_g17255 ( .A(I23341), .ZN(g17255) );
INV_X32 U_g17258 ( .A(g16053), .ZN(g17258) );
INV_X32 U_I23345 ( .A(g15723), .ZN(I23345) );
INV_X32 U_g17259 ( .A(I23345), .ZN(g17259) );
INV_X32 U_I23348 ( .A(g15786), .ZN(I23348) );
INV_X32 U_g17262 ( .A(I23348), .ZN(g17262) );
INV_X32 U_I23351 ( .A(g15788), .ZN(I23351) );
INV_X32 U_g17265 ( .A(I23351), .ZN(g17265) );
INV_X32 U_I23358 ( .A(g16442), .ZN(I23358) );
INV_X32 U_g17272 ( .A(I23358), .ZN(g17272) );
INV_X32 U_I23361 ( .A(g15759), .ZN(I23361) );
INV_X32 U_g17275 ( .A(I23361), .ZN(g17275) );
INV_X32 U_I23364 ( .A(g15805), .ZN(I23364) );
INV_X32 U_g17278 ( .A(I23364), .ZN(g17278) );
INV_X32 U_g17281 ( .A(g16081), .ZN(g17281) );
INV_X32 U_I23368 ( .A(g16446), .ZN(I23368) );
INV_X32 U_g17282 ( .A(I23368), .ZN(g17282) );
INV_X32 U_I23371 ( .A(g15761), .ZN(I23371) );
INV_X32 U_g17285 ( .A(I23371), .ZN(g17285) );
INV_X32 U_I23374 ( .A(g15807), .ZN(I23374) );
INV_X32 U_g17288 ( .A(I23374), .ZN(g17288) );
INV_X32 U_I23377 ( .A(g15763), .ZN(I23377) );
INV_X32 U_g17291 ( .A(I23377), .ZN(g17291) );
INV_X32 U_I23380 ( .A(g15809), .ZN(I23380) );
INV_X32 U_g17294 ( .A(I23380), .ZN(g17294) );
INV_X32 U_I23383 ( .A(g15811), .ZN(I23383) );
INV_X32 U_g17297 ( .A(I23383), .ZN(g17297) );
INV_X32 U_I23386 ( .A(g13469), .ZN(I23386) );
INV_X32 U_g17300 ( .A(I23386), .ZN(g17300) );
INV_X32 U_I23392 ( .A(g13476), .ZN(I23392) );
INV_X32 U_g17304 ( .A(I23392), .ZN(g17304) );
INV_X32 U_I23395 ( .A(g15785), .ZN(I23395) );
INV_X32 U_g17307 ( .A(I23395), .ZN(g17307) );
INV_X32 U_I23398 ( .A(g15820), .ZN(I23398) );
INV_X32 U_g17310 ( .A(I23398), .ZN(g17310) );
INV_X32 U_g17313 ( .A(g16109), .ZN(g17313) );
INV_X32 U_g17314 ( .A(g16110), .ZN(g17314) );
INV_X32 U_I23403 ( .A(g13478), .ZN(I23403) );
INV_X32 U_g17315 ( .A(I23403), .ZN(g17315) );
INV_X32 U_I23406 ( .A(g15787), .ZN(I23406) );
INV_X32 U_g17318 ( .A(I23406), .ZN(g17318) );
INV_X32 U_I23409 ( .A(g15822), .ZN(I23409) );
INV_X32 U_g17321 ( .A(I23409), .ZN(g17321) );
INV_X32 U_I23412 ( .A(g13482), .ZN(I23412) );
INV_X32 U_g17324 ( .A(I23412), .ZN(g17324) );
INV_X32 U_I23415 ( .A(g15789), .ZN(I23415) );
INV_X32 U_g17327 ( .A(I23415), .ZN(g17327) );
INV_X32 U_I23418 ( .A(g15824), .ZN(I23418) );
INV_X32 U_g17330 ( .A(I23418), .ZN(g17330) );
INV_X32 U_I23421 ( .A(g15791), .ZN(I23421) );
INV_X32 U_g17333 ( .A(I23421), .ZN(g17333) );
INV_X32 U_I23424 ( .A(g15826), .ZN(I23424) );
INV_X32 U_g17336 ( .A(I23424), .ZN(g17336) );
INV_X32 U_I23430 ( .A(g13494), .ZN(I23430) );
INV_X32 U_g17342 ( .A(I23430), .ZN(g17342) );
INV_X32 U_I23433 ( .A(g15806), .ZN(I23433) );
INV_X32 U_g17345 ( .A(I23433), .ZN(g17345) );
INV_X32 U_I23436 ( .A(g15832), .ZN(I23436) );
INV_X32 U_g17348 ( .A(I23436), .ZN(g17348) );
INV_X32 U_g17351 ( .A(g16152), .ZN(g17351) );
INV_X32 U_I23442 ( .A(g13495), .ZN(I23442) );
INV_X32 U_g17354 ( .A(I23442), .ZN(g17354) );
INV_X32 U_I23445 ( .A(g15808), .ZN(I23445) );
INV_X32 U_g17357 ( .A(I23445), .ZN(g17357) );
INV_X32 U_I23448 ( .A(g15834), .ZN(I23448) );
INV_X32 U_g17360 ( .A(I23448), .ZN(g17360) );
INV_X32 U_I23451 ( .A(g13497), .ZN(I23451) );
INV_X32 U_g17363 ( .A(I23451), .ZN(g17363) );
INV_X32 U_I23454 ( .A(g15810), .ZN(I23454) );
INV_X32 U_g17366 ( .A(I23454), .ZN(g17366) );
INV_X32 U_I23457 ( .A(g15836), .ZN(I23457) );
INV_X32 U_g17369 ( .A(I23457), .ZN(g17369) );
INV_X32 U_I23460 ( .A(g13501), .ZN(I23460) );
INV_X32 U_g17372 ( .A(I23460), .ZN(g17372) );
INV_X32 U_I23463 ( .A(g15812), .ZN(I23463) );
INV_X32 U_g17375 ( .A(I23463), .ZN(g17375) );
INV_X32 U_I23466 ( .A(g15838), .ZN(I23466) );
INV_X32 U_g17378 ( .A(I23466), .ZN(g17378) );
INV_X32 U_I23472 ( .A(g13510), .ZN(I23472) );
INV_X32 U_g17384 ( .A(I23472), .ZN(g17384) );
INV_X32 U_I23475 ( .A(g15821), .ZN(I23475) );
INV_X32 U_g17387 ( .A(I23475), .ZN(g17387) );
INV_X32 U_I23478 ( .A(g15844), .ZN(I23478) );
INV_X32 U_g17390 ( .A(I23478), .ZN(g17390) );
INV_X32 U_g17394 ( .A(g16197), .ZN(g17394) );
INV_X32 U_I23487 ( .A(g13511), .ZN(I23487) );
INV_X32 U_g17399 ( .A(I23487), .ZN(g17399) );
INV_X32 U_I23490 ( .A(g15823), .ZN(I23490) );
INV_X32 U_g17402 ( .A(I23490), .ZN(g17402) );
INV_X32 U_I23493 ( .A(g15846), .ZN(I23493) );
INV_X32 U_g17405 ( .A(I23493), .ZN(g17405) );
INV_X32 U_I23498 ( .A(g13512), .ZN(I23498) );
INV_X32 U_g17410 ( .A(I23498), .ZN(g17410) );
INV_X32 U_I23501 ( .A(g15825), .ZN(I23501) );
INV_X32 U_g17413 ( .A(I23501), .ZN(g17413) );
INV_X32 U_I23504 ( .A(g15848), .ZN(I23504) );
INV_X32 U_g17416 ( .A(I23504), .ZN(g17416) );
INV_X32 U_I23507 ( .A(g13514), .ZN(I23507) );
INV_X32 U_g17419 ( .A(I23507), .ZN(g17419) );
INV_X32 U_I23510 ( .A(g15827), .ZN(I23510) );
INV_X32 U_g17422 ( .A(I23510), .ZN(g17422) );
INV_X32 U_I23513 ( .A(g15850), .ZN(I23513) );
INV_X32 U_g17425 ( .A(I23513), .ZN(g17425) );
INV_X32 U_I23518 ( .A(g15856), .ZN(I23518) );
INV_X32 U_g17430 ( .A(I23518), .ZN(g17430) );
INV_X32 U_I23521 ( .A(g13518), .ZN(I23521) );
INV_X32 U_g17433 ( .A(I23521), .ZN(g17433) );
INV_X32 U_I23524 ( .A(g15833), .ZN(I23524) );
INV_X32 U_g17436 ( .A(I23524), .ZN(g17436) );
INV_X32 U_I23527 ( .A(g15858), .ZN(I23527) );
INV_X32 U_g17439 ( .A(I23527), .ZN(g17439) );
INV_X32 U_I23530 ( .A(g14885), .ZN(I23530) );
INV_X32 U_g17442 ( .A(I23530), .ZN(g17442) );
INV_X32 U_g17445 ( .A(g16250), .ZN(g17445) );
INV_X32 U_I23539 ( .A(g13524), .ZN(I23539) );
INV_X32 U_g17451 ( .A(I23539), .ZN(g17451) );
INV_X32 U_I23542 ( .A(g15835), .ZN(I23542) );
INV_X32 U_g17454 ( .A(I23542), .ZN(g17454) );
INV_X32 U_I23545 ( .A(g15867), .ZN(I23545) );
INV_X32 U_g17457 ( .A(I23545), .ZN(g17457) );
INV_X32 U_I23553 ( .A(g13525), .ZN(I23553) );
INV_X32 U_g17465 ( .A(I23553), .ZN(g17465) );
INV_X32 U_I23556 ( .A(g15837), .ZN(I23556) );
INV_X32 U_g17468 ( .A(I23556), .ZN(g17468) );
INV_X32 U_I23559 ( .A(g15869), .ZN(I23559) );
INV_X32 U_g17471 ( .A(I23559), .ZN(g17471) );
INV_X32 U_I23564 ( .A(g13526), .ZN(I23564) );
INV_X32 U_g17476 ( .A(I23564), .ZN(g17476) );
INV_X32 U_I23567 ( .A(g15839), .ZN(I23567) );
INV_X32 U_g17479 ( .A(I23567), .ZN(g17479) );
INV_X32 U_I23570 ( .A(g15871), .ZN(I23570) );
INV_X32 U_g17482 ( .A(I23570), .ZN(g17482) );
INV_X32 U_I23575 ( .A(g15843), .ZN(I23575) );
INV_X32 U_g17487 ( .A(I23575), .ZN(g17487) );
INV_X32 U_I23578 ( .A(g15879), .ZN(I23578) );
INV_X32 U_g17490 ( .A(I23578), .ZN(g17490) );
INV_X32 U_I23581 ( .A(g13528), .ZN(I23581) );
INV_X32 U_g17493 ( .A(I23581), .ZN(g17493) );
INV_X32 U_I23584 ( .A(g15845), .ZN(I23584) );
INV_X32 U_g17496 ( .A(I23584), .ZN(g17496) );
INV_X32 U_g17499 ( .A(g16292), .ZN(g17499) );
INV_X32 U_I23588 ( .A(g14885), .ZN(I23588) );
INV_X32 U_g17500 ( .A(I23588), .ZN(g17500) );
INV_X32 U_I23591 ( .A(g14885), .ZN(I23591) );
INV_X32 U_g17503 ( .A(I23591), .ZN(g17503) );
INV_X32 U_I23599 ( .A(g15887), .ZN(I23599) );
INV_X32 U_g17511 ( .A(I23599), .ZN(g17511) );
INV_X32 U_I23602 ( .A(g13529), .ZN(I23602) );
INV_X32 U_g17514 ( .A(I23602), .ZN(g17514) );
INV_X32 U_I23605 ( .A(g15847), .ZN(I23605) );
INV_X32 U_g17517 ( .A(I23605), .ZN(g17517) );
INV_X32 U_I23608 ( .A(g15889), .ZN(I23608) );
INV_X32 U_g17520 ( .A(I23608), .ZN(g17520) );
INV_X32 U_I23611 ( .A(g14966), .ZN(I23611) );
INV_X32 U_g17523 ( .A(I23611), .ZN(g17523) );
INV_X32 U_I23619 ( .A(g13535), .ZN(I23619) );
INV_X32 U_g17531 ( .A(I23619), .ZN(g17531) );
INV_X32 U_I23622 ( .A(g15849), .ZN(I23622) );
INV_X32 U_g17534 ( .A(I23622), .ZN(g17534) );
INV_X32 U_I23625 ( .A(g15898), .ZN(I23625) );
INV_X32 U_g17537 ( .A(I23625), .ZN(g17537) );
INV_X32 U_I23633 ( .A(g13536), .ZN(I23633) );
INV_X32 U_g17545 ( .A(I23633), .ZN(g17545) );
INV_X32 U_I23636 ( .A(g15851), .ZN(I23636) );
INV_X32 U_g17548 ( .A(I23636), .ZN(g17548) );
INV_X32 U_I23639 ( .A(g15900), .ZN(I23639) );
INV_X32 U_g17551 ( .A(I23639), .ZN(g17551) );
INV_X32 U_I23645 ( .A(g13537), .ZN(I23645) );
INV_X32 U_g17557 ( .A(I23645), .ZN(g17557) );
INV_X32 U_I23648 ( .A(g15857), .ZN(I23648) );
INV_X32 U_g17560 ( .A(I23648), .ZN(g17560) );
INV_X32 U_I23651 ( .A(g13538), .ZN(I23651) );
INV_X32 U_g17563 ( .A(I23651), .ZN(g17563) );
INV_X32 U_g17566 ( .A(g16346), .ZN(g17566) );
INV_X32 U_I23655 ( .A(g14831), .ZN(I23655) );
INV_X32 U_g17567 ( .A(I23655), .ZN(g17567) );
INV_X32 U_I23658 ( .A(g14885), .ZN(I23658) );
INV_X32 U_g17570 ( .A(I23658), .ZN(g17570) );
INV_X32 U_I23661 ( .A(g16085), .ZN(I23661) );
INV_X32 U_g17573 ( .A(I23661), .ZN(g17573) );
INV_X32 U_I23667 ( .A(g15866), .ZN(I23667) );
INV_X32 U_g17579 ( .A(I23667), .ZN(g17579) );
INV_X32 U_I23670 ( .A(g15912), .ZN(I23670) );
INV_X32 U_g17582 ( .A(I23670), .ZN(g17582) );
INV_X32 U_I23673 ( .A(g13539), .ZN(I23673) );
INV_X32 U_g17585 ( .A(I23673), .ZN(g17585) );
INV_X32 U_I23676 ( .A(g15868), .ZN(I23676) );
INV_X32 U_g17588 ( .A(I23676), .ZN(g17588) );
INV_X32 U_I23679 ( .A(g14966), .ZN(I23679) );
INV_X32 U_g17591 ( .A(I23679), .ZN(g17591) );
INV_X32 U_I23682 ( .A(g14966), .ZN(I23682) );
INV_X32 U_g17594 ( .A(I23682), .ZN(g17594) );
INV_X32 U_I23689 ( .A(g15920), .ZN(I23689) );
INV_X32 U_g17601 ( .A(I23689), .ZN(g17601) );
INV_X32 U_I23692 ( .A(g13540), .ZN(I23692) );
INV_X32 U_g17604 ( .A(I23692), .ZN(g17604) );
INV_X32 U_I23695 ( .A(g15870), .ZN(I23695) );
INV_X32 U_g17607 ( .A(I23695), .ZN(g17607) );
INV_X32 U_I23698 ( .A(g15922), .ZN(I23698) );
INV_X32 U_g17610 ( .A(I23698), .ZN(g17610) );
INV_X32 U_I23701 ( .A(g15055), .ZN(I23701) );
INV_X32 U_g17613 ( .A(I23701), .ZN(g17613) );
INV_X32 U_I23709 ( .A(g13546), .ZN(I23709) );
INV_X32 U_g17621 ( .A(I23709), .ZN(g17621) );
INV_X32 U_I23712 ( .A(g15872), .ZN(I23712) );
INV_X32 U_g17624 ( .A(I23712), .ZN(g17624) );
INV_X32 U_I23715 ( .A(g15931), .ZN(I23715) );
INV_X32 U_g17627 ( .A(I23715), .ZN(g17627) );
INV_X32 U_I23725 ( .A(g13547), .ZN(I23725) );
INV_X32 U_g17637 ( .A(I23725), .ZN(g17637) );
INV_X32 U_g17640 ( .A(g13873), .ZN(g17640) );
INV_X32 U_I23729 ( .A(g14337), .ZN(I23729) );
INV_X32 U_g17645 ( .A(I23729), .ZN(g17645) );
INV_X32 U_g17648 ( .A(g16384), .ZN(g17648) );
INV_X32 U_I23733 ( .A(g14831), .ZN(I23733) );
INV_X32 U_g17649 ( .A(I23733), .ZN(g17649) );
INV_X32 U_I23739 ( .A(g13548), .ZN(I23739) );
INV_X32 U_g17655 ( .A(I23739), .ZN(g17655) );
INV_X32 U_I23742 ( .A(g15888), .ZN(I23742) );
INV_X32 U_g17658 ( .A(I23742), .ZN(g17658) );
INV_X32 U_I23745 ( .A(g13549), .ZN(I23745) );
INV_X32 U_g17661 ( .A(I23745), .ZN(g17661) );
INV_X32 U_I23748 ( .A(g14904), .ZN(I23748) );
INV_X32 U_g17664 ( .A(I23748), .ZN(g17664) );
INV_X32 U_I23751 ( .A(g14966), .ZN(I23751) );
INV_X32 U_g17667 ( .A(I23751), .ZN(g17667) );
INV_X32 U_I23754 ( .A(g16123), .ZN(I23754) );
INV_X32 U_g17670 ( .A(I23754), .ZN(g17670) );
INV_X32 U_I23760 ( .A(g15897), .ZN(I23760) );
INV_X32 U_g17676 ( .A(I23760), .ZN(g17676) );
INV_X32 U_I23763 ( .A(g15941), .ZN(I23763) );
INV_X32 U_g17679 ( .A(I23763), .ZN(g17679) );
INV_X32 U_I23766 ( .A(g13550), .ZN(I23766) );
INV_X32 U_g17682 ( .A(I23766), .ZN(g17682) );
INV_X32 U_I23769 ( .A(g15899), .ZN(I23769) );
INV_X32 U_g17685 ( .A(I23769), .ZN(g17685) );
INV_X32 U_I23772 ( .A(g15055), .ZN(I23772) );
INV_X32 U_g17688 ( .A(I23772), .ZN(g17688) );
INV_X32 U_I23775 ( .A(g15055), .ZN(I23775) );
INV_X32 U_g17691 ( .A(I23775), .ZN(g17691) );
INV_X32 U_I23782 ( .A(g15949), .ZN(I23782) );
INV_X32 U_g17698 ( .A(I23782), .ZN(g17698) );
INV_X32 U_I23785 ( .A(g13551), .ZN(I23785) );
INV_X32 U_g17701 ( .A(I23785), .ZN(g17701) );
INV_X32 U_I23788 ( .A(g15901), .ZN(I23788) );
INV_X32 U_g17704 ( .A(I23788), .ZN(g17704) );
INV_X32 U_I23791 ( .A(g15951), .ZN(I23791) );
INV_X32 U_g17707 ( .A(I23791), .ZN(g17707) );
INV_X32 U_I23794 ( .A(g15151), .ZN(I23794) );
INV_X32 U_g17710 ( .A(I23794), .ZN(g17710) );
INV_X32 U_g17720 ( .A(g15853), .ZN(g17720) );
INV_X32 U_g17724 ( .A(g13886), .ZN(g17724) );
INV_X32 U_I23817 ( .A(g13557), .ZN(I23817) );
INV_X32 U_g17738 ( .A(I23817), .ZN(g17738) );
INV_X32 U_g17741 ( .A(g13895), .ZN(g17741) );
INV_X32 U_I23821 ( .A(g14337), .ZN(I23821) );
INV_X32 U_g17746 ( .A(I23821), .ZN(g17746) );
INV_X32 U_I23824 ( .A(g14904), .ZN(I23824) );
INV_X32 U_g17749 ( .A(I23824), .ZN(g17749) );
INV_X32 U_I23830 ( .A(g13558), .ZN(I23830) );
INV_X32 U_g17755 ( .A(I23830), .ZN(g17755) );
INV_X32 U_I23833 ( .A(g15921), .ZN(I23833) );
INV_X32 U_g17758 ( .A(I23833), .ZN(g17758) );
INV_X32 U_I23836 ( .A(g13559), .ZN(I23836) );
INV_X32 U_g17761 ( .A(I23836), .ZN(g17761) );
INV_X32 U_I23839 ( .A(g14985), .ZN(I23839) );
INV_X32 U_g17764 ( .A(I23839), .ZN(g17764) );
INV_X32 U_I23842 ( .A(g15055), .ZN(I23842) );
INV_X32 U_g17767 ( .A(I23842), .ZN(g17767) );
INV_X32 U_I23845 ( .A(g16174), .ZN(I23845) );
INV_X32 U_g17770 ( .A(I23845), .ZN(g17770) );
INV_X32 U_I23851 ( .A(g15930), .ZN(I23851) );
INV_X32 U_g17776 ( .A(I23851), .ZN(g17776) );
INV_X32 U_I23854 ( .A(g15970), .ZN(I23854) );
INV_X32 U_g17779 ( .A(I23854), .ZN(g17779) );
INV_X32 U_I23857 ( .A(g13560), .ZN(I23857) );
INV_X32 U_g17782 ( .A(I23857), .ZN(g17782) );
INV_X32 U_I23860 ( .A(g15932), .ZN(I23860) );
INV_X32 U_g17785 ( .A(I23860), .ZN(g17785) );
INV_X32 U_I23863 ( .A(g15151), .ZN(I23863) );
INV_X32 U_g17788 ( .A(I23863), .ZN(g17788) );
INV_X32 U_I23866 ( .A(g15151), .ZN(I23866) );
INV_X32 U_g17791 ( .A(I23866), .ZN(g17791) );
INV_X32 U_I23874 ( .A(g15797), .ZN(I23874) );
INV_X32 U_g17799 ( .A(I23874), .ZN(g17799) );
INV_X32 U_g17802 ( .A(g13907), .ZN(g17802) );
INV_X32 U_I23888 ( .A(g14685), .ZN(I23888) );
INV_X32 U_g17815 ( .A(I23888), .ZN(g17815) );
INV_X32 U_g17825 ( .A(g13927), .ZN(g17825) );
INV_X32 U_I23904 ( .A(g13561), .ZN(I23904) );
INV_X32 U_g17839 ( .A(I23904), .ZN(g17839) );
INV_X32 U_g17842 ( .A(g13936), .ZN(g17842) );
INV_X32 U_I23908 ( .A(g14337), .ZN(I23908) );
INV_X32 U_g17847 ( .A(I23908), .ZN(g17847) );
INV_X32 U_I23911 ( .A(g14985), .ZN(I23911) );
INV_X32 U_g17850 ( .A(I23911), .ZN(g17850) );
INV_X32 U_I23917 ( .A(g13562), .ZN(I23917) );
INV_X32 U_g17856 ( .A(I23917), .ZN(g17856) );
INV_X32 U_I23920 ( .A(g15950), .ZN(I23920) );
INV_X32 U_g17859 ( .A(I23920), .ZN(g17859) );
INV_X32 U_I23923 ( .A(g13563), .ZN(I23923) );
INV_X32 U_g17862 ( .A(I23923), .ZN(g17862) );
INV_X32 U_I23926 ( .A(g15074), .ZN(I23926) );
INV_X32 U_g17865 ( .A(I23926), .ZN(g17865) );
INV_X32 U_I23929 ( .A(g15151), .ZN(I23929) );
INV_X32 U_g17868 ( .A(I23929), .ZN(g17868) );
INV_X32 U_I23932 ( .A(g16233), .ZN(I23932) );
INV_X32 U_g17871 ( .A(I23932), .ZN(g17871) );
INV_X32 U_g17878 ( .A(g15830), .ZN(g17878) );
INV_X32 U_g17882 ( .A(g13946), .ZN(g17882) );
INV_X32 U_g17892 ( .A(g13954), .ZN(g17892) );
INV_X32 U_g17893 ( .A(g14165), .ZN(g17893) );
INV_X32 U_I23954 ( .A(g16154), .ZN(I23954) );
INV_X32 U_g17903 ( .A(I23954), .ZN(g17903) );
INV_X32 U_g17914 ( .A(g13963), .ZN(g17914) );
INV_X32 U_I23976 ( .A(g14719), .ZN(I23976) );
INV_X32 U_g17927 ( .A(I23976), .ZN(g17927) );
INV_X32 U_g17937 ( .A(g13983), .ZN(g17937) );
INV_X32 U_I23992 ( .A(g13564), .ZN(I23992) );
INV_X32 U_g17951 ( .A(I23992), .ZN(g17951) );
INV_X32 U_g17954 ( .A(g13992), .ZN(g17954) );
INV_X32 U_I23996 ( .A(g14337), .ZN(I23996) );
INV_X32 U_g17959 ( .A(I23996), .ZN(g17959) );
INV_X32 U_I23999 ( .A(g15074), .ZN(I23999) );
INV_X32 U_g17962 ( .A(I23999), .ZN(g17962) );
INV_X32 U_g17969 ( .A(g15841), .ZN(g17969) );
INV_X32 U_g17974 ( .A(g14001), .ZN(g17974) );
INV_X32 U_g17984 ( .A(g14008), .ZN(g17984) );
INV_X32 U_g17988 ( .A(g14685), .ZN(g17988) );
INV_X32 U_g17991 ( .A(g14450), .ZN(g17991) );
INV_X32 U_g17993 ( .A(g14016), .ZN(g17993) );
INV_X32 U_g18003 ( .A(g14024), .ZN(g18003) );
INV_X32 U_g18004 ( .A(g14280), .ZN(g18004) );
INV_X32 U_I24049 ( .A(g16213), .ZN(I24049) );
INV_X32 U_g18014 ( .A(I24049), .ZN(g18014) );
INV_X32 U_g18025 ( .A(g14033), .ZN(g18025) );
INV_X32 U_I24071 ( .A(g14747), .ZN(I24071) );
INV_X32 U_g18038 ( .A(I24071), .ZN(g18038) );
INV_X32 U_g18048 ( .A(g14053), .ZN(g18048) );
INV_X32 U_g18063 ( .A(g15660), .ZN(g18063) );
INV_X32 U_g18070 ( .A(g15854), .ZN(g18070) );
INV_X32 U_g18074 ( .A(g14062), .ZN(g18074) );
INV_X32 U_g18084 ( .A(g14068), .ZN(g18084) );
INV_X32 U_g18089 ( .A(g14355), .ZN(g18089) );
INV_X32 U_g18091 ( .A(g14092), .ZN(g18091) );
INV_X32 U_g18101 ( .A(g14099), .ZN(g18101) );
INV_X32 U_g18105 ( .A(g14719), .ZN(g18105) );
INV_X32 U_g18108 ( .A(g14537), .ZN(g18108) );
INV_X32 U_g18110 ( .A(g14107), .ZN(g18110) );
INV_X32 U_g18120 ( .A(g14115), .ZN(g18120) );
INV_X32 U_g18121 ( .A(g14402), .ZN(g18121) );
INV_X32 U_I24144 ( .A(g16278), .ZN(I24144) );
INV_X32 U_g18131 ( .A(I24144), .ZN(g18131) );
INV_X32 U_g18142 ( .A(g14124), .ZN(g18142) );
INV_X32 U_I24166 ( .A(g14768), .ZN(I24166) );
INV_X32 U_g18155 ( .A(I24166), .ZN(g18155) );
INV_X32 U_I24171 ( .A(g16439), .ZN(I24171) );
INV_X32 U_g18166 ( .A(I24171), .ZN(g18166) );
INV_X32 U_g18170 ( .A(g15877), .ZN(g18170) );
INV_X32 U_g18174 ( .A(g14148), .ZN(g18174) );
INV_X32 U_g18179 ( .A(g14153), .ZN(g18179) );
INV_X32 U_g18188 ( .A(g14252), .ZN(g18188) );
INV_X32 U_g18190 ( .A(g14177), .ZN(g18190) );
INV_X32 U_g18200 ( .A(g14183), .ZN(g18200) );
INV_X32 U_g18205 ( .A(g14467), .ZN(g18205) );
INV_X32 U_g18207 ( .A(g14207), .ZN(g18207) );
INV_X32 U_g18217 ( .A(g14214), .ZN(g18217) );
INV_X32 U_g18221 ( .A(g14747), .ZN(g18221) );
INV_X32 U_g18224 ( .A(g14592), .ZN(g18224) );
INV_X32 U_g18226 ( .A(g14222), .ZN(g18226) );
INV_X32 U_g18236 ( .A(g14230), .ZN(g18236) );
INV_X32 U_g18237 ( .A(g14514), .ZN(g18237) );
INV_X32 U_I24247 ( .A(g16337), .ZN(I24247) );
INV_X32 U_g18247 ( .A(I24247), .ZN(g18247) );
INV_X32 U_I24258 ( .A(g16463), .ZN(I24258) );
INV_X32 U_g18258 ( .A(I24258), .ZN(g18258) );
INV_X32 U_g18261 ( .A(g15719), .ZN(g18261) );
INV_X32 U_g18265 ( .A(g14238), .ZN(g18265) );
INV_X32 U_g18275 ( .A(g14171), .ZN(g18275) );
INV_X32 U_I24285 ( .A(g15992), .ZN(I24285) );
INV_X32 U_g18278 ( .A(I24285), .ZN(g18278) );
INV_X32 U_g18281 ( .A(g14263), .ZN(g18281) );
INV_X32 U_g18286 ( .A(g14268), .ZN(g18286) );
INV_X32 U_g18295 ( .A(g14374), .ZN(g18295) );
INV_X32 U_g18297 ( .A(g14292), .ZN(g18297) );
INV_X32 U_g18307 ( .A(g14298), .ZN(g18307) );
INV_X32 U_g18312 ( .A(g14554), .ZN(g18312) );
INV_X32 U_g18314 ( .A(g14322), .ZN(g18314) );
INV_X32 U_g18324 ( .A(g14329), .ZN(g18324) );
INV_X32 U_g18328 ( .A(g14768), .ZN(g18328) );
INV_X32 U_g18331 ( .A(g14626), .ZN(g18331) );
INV_X32 U_I24346 ( .A(g15873), .ZN(I24346) );
INV_X32 U_g18334 ( .A(I24346), .ZN(g18334) );
INV_X32 U_g18337 ( .A(g15757), .ZN(g18337) );
INV_X32 U_g18341 ( .A(g14342), .ZN(g18341) );
INV_X32 U_g18351 ( .A(g13741), .ZN(g18351) );
INV_X32 U_g18353 ( .A(g13918), .ZN(g18353) );
INV_X32 U_I24368 ( .A(g15990), .ZN(I24368) );
INV_X32 U_g18355 ( .A(I24368), .ZN(g18355) );
INV_X32 U_g18358 ( .A(g14360), .ZN(g18358) );
INV_X32 U_g18368 ( .A(g14286), .ZN(g18368) );
INV_X32 U_I24394 ( .A(g15995), .ZN(I24394) );
INV_X32 U_g18371 ( .A(I24394), .ZN(g18371) );
INV_X32 U_g18374 ( .A(g14385), .ZN(g18374) );
INV_X32 U_g18379 ( .A(g14390), .ZN(g18379) );
INV_X32 U_g18388 ( .A(g14486), .ZN(g18388) );
INV_X32 U_g18390 ( .A(g14414), .ZN(g18390) );
INV_X32 U_g18400 ( .A(g14420), .ZN(g18400) );
INV_X32 U_g18405 ( .A(g14609), .ZN(g18405) );
INV_X32 U_g18407 ( .A(g15959), .ZN(g18407) );
INV_X32 U_g18414 ( .A(g15718), .ZN(g18414) );
INV_X32 U_g18415 ( .A(g15783), .ZN(g18415) );
INV_X32 U_g18429 ( .A(g14831), .ZN(g18429) );
INV_X32 U_I24459 ( .A(g13599), .ZN(I24459) );
INV_X32 U_g18432 ( .A(I24459), .ZN(g18432) );
INV_X32 U_g18435 ( .A(g14359), .ZN(g18435) );
INV_X32 U_g18436 ( .A(g14454), .ZN(g18436) );
INV_X32 U_g18446 ( .A(g13741), .ZN(g18446) );
INV_X32 U_g18448 ( .A(g13974), .ZN(g18448) );
INV_X32 U_I24481 ( .A(g15993), .ZN(I24481) );
INV_X32 U_g18450 ( .A(I24481), .ZN(g18450) );
INV_X32 U_g18453 ( .A(g14472), .ZN(g18453) );
INV_X32 U_g18463 ( .A(g14408), .ZN(g18463) );
INV_X32 U_I24507 ( .A(g15999), .ZN(I24507) );
INV_X32 U_g18466 ( .A(I24507), .ZN(g18466) );
INV_X32 U_g18469 ( .A(g14497), .ZN(g18469) );
INV_X32 U_g18474 ( .A(g14502), .ZN(g18474) );
INV_X32 U_g18483 ( .A(g14573), .ZN(g18483) );
INV_X32 U_g18485 ( .A(g15756), .ZN(g18485) );
INV_X32 U_g18486 ( .A(g15804), .ZN(g18486) );
INV_X32 U_g18490 ( .A(g13565), .ZN(g18490) );
INV_X32 U_g18502 ( .A(g14904), .ZN(g18502) );
INV_X32 U_I24560 ( .A(g13611), .ZN(I24560) );
INV_X32 U_g18505 ( .A(I24560), .ZN(g18505) );
INV_X32 U_g18508 ( .A(g14471), .ZN(g18508) );
INV_X32 U_g18509 ( .A(g14541), .ZN(g18509) );
INV_X32 U_g18519 ( .A(g13741), .ZN(g18519) );
INV_X32 U_g18521 ( .A(g14044), .ZN(g18521) );
INV_X32 U_I24582 ( .A(g15996), .ZN(I24582) );
INV_X32 U_g18523 ( .A(I24582), .ZN(g18523) );
INV_X32 U_g18526 ( .A(g14559), .ZN(g18526) );
INV_X32 U_g18536 ( .A(g14520), .ZN(g18536) );
INV_X32 U_I24608 ( .A(g16006), .ZN(I24608) );
INV_X32 U_g18539 ( .A(I24608), .ZN(g18539) );
INV_X32 U_g18543 ( .A(g15819), .ZN(g18543) );
INV_X32 U_g18552 ( .A(g16154), .ZN(g18552) );
INV_X32 U_g18554 ( .A(g13573), .ZN(g18554) );
INV_X32 U_g18566 ( .A(g14985), .ZN(g18566) );
INV_X32 U_I24662 ( .A(g13621), .ZN(I24662) );
INV_X32 U_g18569 ( .A(I24662), .ZN(g18569) );
INV_X32 U_g18572 ( .A(g14558), .ZN(g18572) );
INV_X32 U_g18573 ( .A(g14596), .ZN(g18573) );
INV_X32 U_g18583 ( .A(g13741), .ZN(g18583) );
INV_X32 U_g18585 ( .A(g14135), .ZN(g18585) );
INV_X32 U_I24684 ( .A(g16000), .ZN(I24684) );
INV_X32 U_g18587 ( .A(I24684), .ZN(g18587) );
INV_X32 U_g18593 ( .A(g15831), .ZN(g18593) );
INV_X32 U_g18602 ( .A(g16213), .ZN(g18602) );
INV_X32 U_g18604 ( .A(g13582), .ZN(g18604) );
INV_X32 U_g18616 ( .A(g15074), .ZN(g18616) );
INV_X32 U_I24732 ( .A(g13633), .ZN(I24732) );
INV_X32 U_g18619 ( .A(I24732), .ZN(g18619) );
INV_X32 U_g18622 ( .A(g14613), .ZN(g18622) );
INV_X32 U_g18634 ( .A(g16278), .ZN(g18634) );
INV_X32 U_g18636 ( .A(g13602), .ZN(g18636) );
INV_X32 U_g18643 ( .A(g16337), .ZN(g18643) );
INV_X32 U_g18646 ( .A(g16341), .ZN(g18646) );
INV_X32 U_g18656 ( .A(g14776), .ZN(g18656) );
INV_X32 U_g18670 ( .A(g14797), .ZN(g18670) );
INV_X32 U_g18679 ( .A(g14811), .ZN(g18679) );
INV_X32 U_g18691 ( .A(g14885), .ZN(g18691) );
INV_X32 U_g18692 ( .A(g14837), .ZN(g18692) );
INV_X32 U_g18699 ( .A(g14849), .ZN(g18699) );
INV_X32 U_g18708 ( .A(g14863), .ZN(g18708) );
INV_X32 U_g18720 ( .A(g14895), .ZN(g18720) );
INV_X32 U_g18725 ( .A(g13865), .ZN(g18725) );
INV_X32 U_g18727 ( .A(g14966), .ZN(g18727) );
INV_X32 U_g18728 ( .A(g14910), .ZN(g18728) );
INV_X32 U_g18735 ( .A(g14922), .ZN(g18735) );
INV_X32 U_g18744 ( .A(g14936), .ZN(g18744) );
INV_X32 U_g18756 ( .A(g14960), .ZN(g18756) );
INV_X32 U_g18757 ( .A(g14963), .ZN(g18757) );
INV_X32 U_g18758 ( .A(g14976), .ZN(g18758) );
INV_X32 U_g18764 ( .A(g15055), .ZN(g18764) );
INV_X32 U_g18765 ( .A(g14991), .ZN(g18765) );
INV_X32 U_g18772 ( .A(g15003), .ZN(g18772) );
INV_X32 U_g18783 ( .A(g15034), .ZN(g18783) );
INV_X32 U_g18784 ( .A(g15037), .ZN(g18784) );
INV_X32 U_g18785 ( .A(g15040), .ZN(g18785) );
INV_X32 U_g18786 ( .A(g15043), .ZN(g18786) );
INV_X32 U_g18787 ( .A(g15049), .ZN(g18787) );
INV_X32 U_g18788 ( .A(g15052), .ZN(g18788) );
INV_X32 U_g18789 ( .A(g15065), .ZN(g18789) );
INV_X32 U_g18795 ( .A(g15151), .ZN(g18795) );
INV_X32 U_g18796 ( .A(g15080), .ZN(g18796) );
INV_X32 U_g18805 ( .A(g15106), .ZN(g18805) );
INV_X32 U_g18806 ( .A(g15109), .ZN(g18806) );
INV_X32 U_g18807 ( .A(g15112), .ZN(g18807) );
INV_X32 U_g18808 ( .A(g15115), .ZN(g18808) );
INV_X32 U_g18809 ( .A(g15130), .ZN(g18809) );
INV_X32 U_g18810 ( .A(g15133), .ZN(g18810) );
INV_X32 U_g18811 ( .A(g15136), .ZN(g18811) );
INV_X32 U_g18812 ( .A(g15139), .ZN(g18812) );
INV_X32 U_g18813 ( .A(g15145), .ZN(g18813) );
INV_X32 U_g18814 ( .A(g15148), .ZN(g18814) );
INV_X32 U_g18815 ( .A(g15161), .ZN(g18815) );
INV_X32 U_g18822 ( .A(g15179), .ZN(g18822) );
INV_X32 U_g18823 ( .A(g15182), .ZN(g18823) );
INV_X32 U_g18824 ( .A(g15185), .ZN(g18824) );
INV_X32 U_g18825 ( .A(g15198), .ZN(g18825) );
INV_X32 U_g18826 ( .A(g15201), .ZN(g18826) );
INV_X32 U_g18827 ( .A(g15204), .ZN(g18827) );
INV_X32 U_g18828 ( .A(g15207), .ZN(g18828) );
INV_X32 U_g18829 ( .A(g15222), .ZN(g18829) );
INV_X32 U_g18830 ( .A(g15225), .ZN(g18830) );
INV_X32 U_g18831 ( .A(g15228), .ZN(g18831) );
INV_X32 U_g18832 ( .A(g15231), .ZN(g18832) );
INV_X32 U_g18833 ( .A(g15237), .ZN(g18833) );
INV_X32 U_g18834 ( .A(g15240), .ZN(g18834) );
INV_X32 U_g18838 ( .A(g15248), .ZN(g18838) );
INV_X32 U_g18839 ( .A(g15251), .ZN(g18839) );
INV_X32 U_g18840 ( .A(g15254), .ZN(g18840) );
INV_X32 U_g18841 ( .A(g15265), .ZN(g18841) );
INV_X32 U_g18842 ( .A(g15268), .ZN(g18842) );
INV_X32 U_g18843 ( .A(g15271), .ZN(g18843) );
INV_X32 U_g18844 ( .A(g15284), .ZN(g18844) );
INV_X32 U_g18845 ( .A(g15287), .ZN(g18845) );
INV_X32 U_g18846 ( .A(g15290), .ZN(g18846) );
INV_X32 U_g18847 ( .A(g15293), .ZN(g18847) );
INV_X32 U_g18848 ( .A(g15308), .ZN(g18848) );
INV_X32 U_g18849 ( .A(g15311), .ZN(g18849) );
INV_X32 U_g18850 ( .A(g15314), .ZN(g18850) );
INV_X32 U_g18851 ( .A(g15317), .ZN(g18851) );
INV_X32 U_g18853 ( .A(g15326), .ZN(g18853) );
INV_X32 U_g18854 ( .A(g15329), .ZN(g18854) );
INV_X32 U_g18855 ( .A(g15332), .ZN(g18855) );
INV_X32 U_g18856 ( .A(g15340), .ZN(g18856) );
INV_X32 U_g18857 ( .A(g15343), .ZN(g18857) );
INV_X32 U_g18858 ( .A(g15346), .ZN(g18858) );
INV_X32 U_g18859 ( .A(g15357), .ZN(g18859) );
INV_X32 U_g18860 ( .A(g15360), .ZN(g18860) );
INV_X32 U_g18861 ( .A(g15363), .ZN(g18861) );
INV_X32 U_g18862 ( .A(g15376), .ZN(g18862) );
INV_X32 U_g18863 ( .A(g15379), .ZN(g18863) );
INV_X32 U_g18864 ( .A(g15382), .ZN(g18864) );
INV_X32 U_g18865 ( .A(g15385), .ZN(g18865) );
INV_X32 U_I24894 ( .A(g14797), .ZN(I24894) );
INV_X32 U_g18869 ( .A(I24894), .ZN(g18869) );
INV_X32 U_g18870 ( .A(g15393), .ZN(g18870) );
INV_X32 U_g18871 ( .A(g15396), .ZN(g18871) );
INV_X32 U_g18872 ( .A(g15399), .ZN(g18872) );
INV_X32 U_g18873 ( .A(g15404), .ZN(g18873) );
INV_X32 U_g18874 ( .A(g15412), .ZN(g18874) );
INV_X32 U_g18875 ( .A(g15415), .ZN(g18875) );
INV_X32 U_g18876 ( .A(g15418), .ZN(g18876) );
INV_X32 U_g18877 ( .A(g15426), .ZN(g18877) );
INV_X32 U_g18878 ( .A(g15429), .ZN(g18878) );
INV_X32 U_g18879 ( .A(g15432), .ZN(g18879) );
INV_X32 U_g18880 ( .A(g15443), .ZN(g18880) );
INV_X32 U_g18881 ( .A(g15446), .ZN(g18881) );
INV_X32 U_g18882 ( .A(g15449), .ZN(g18882) );
INV_X32 U_g18884 ( .A(g13469), .ZN(g18884) );
INV_X32 U_I24913 ( .A(g15800), .ZN(I24913) );
INV_X32 U_g18886 ( .A(I24913), .ZN(g18886) );
INV_X32 U_I24916 ( .A(g14776), .ZN(I24916) );
INV_X32 U_g18890 ( .A(I24916), .ZN(g18890) );
INV_X32 U_g18891 ( .A(g15461), .ZN(g18891) );
INV_X32 U_g18892 ( .A(g15464), .ZN(g18892) );
INV_X32 U_g18893 ( .A(g15467), .ZN(g18893) );
INV_X32 U_g18894 ( .A(g15471), .ZN(g18894) );
INV_X32 U_I24923 ( .A(g14849), .ZN(I24923) );
INV_X32 U_g18895 ( .A(I24923), .ZN(g18895) );
INV_X32 U_g18896 ( .A(g15477), .ZN(g18896) );
INV_X32 U_g18897 ( .A(g15480), .ZN(g18897) );
INV_X32 U_g18898 ( .A(g15483), .ZN(g18898) );
INV_X32 U_g18899 ( .A(g15488), .ZN(g18899) );
INV_X32 U_g18900 ( .A(g15496), .ZN(g18900) );
INV_X32 U_g18901 ( .A(g15499), .ZN(g18901) );
INV_X32 U_g18902 ( .A(g15502), .ZN(g18902) );
INV_X32 U_g18903 ( .A(g15510), .ZN(g18903) );
INV_X32 U_g18904 ( .A(g15513), .ZN(g18904) );
INV_X32 U_g18905 ( .A(g15516), .ZN(g18905) );
INV_X32 U_g18908 ( .A(g15521), .ZN(g18908) );
INV_X32 U_g18909 ( .A(g15528), .ZN(g18909) );
INV_X32 U_g18910 ( .A(g15531), .ZN(g18910) );
INV_X32 U_g18911 ( .A(g15534), .ZN(g18911) );
INV_X32 U_g18912 ( .A(g15537), .ZN(g18912) );
INV_X32 U_I24943 ( .A(g14811), .ZN(I24943) );
INV_X32 U_g18913 ( .A(I24943), .ZN(g18913) );
INV_X32 U_g18914 ( .A(g15547), .ZN(g18914) );
INV_X32 U_g18915 ( .A(g15550), .ZN(g18915) );
INV_X32 U_g18916 ( .A(g15553), .ZN(g18916) );
INV_X32 U_g18917 ( .A(g15557), .ZN(g18917) );
INV_X32 U_I24950 ( .A(g14922), .ZN(I24950) );
INV_X32 U_g18918 ( .A(I24950), .ZN(g18918) );
INV_X32 U_g18919 ( .A(g15563), .ZN(g18919) );
INV_X32 U_g18920 ( .A(g15566), .ZN(g18920) );
INV_X32 U_g18921 ( .A(g15569), .ZN(g18921) );
INV_X32 U_g18922 ( .A(g15574), .ZN(g18922) );
INV_X32 U_g18923 ( .A(g15582), .ZN(g18923) );
INV_X32 U_g18924 ( .A(g15585), .ZN(g18924) );
INV_X32 U_g18925 ( .A(g15588), .ZN(g18925) );
INV_X32 U_g18926 ( .A(g15596), .ZN(g18926) );
INV_X32 U_g18927 ( .A(g15599), .ZN(g18927) );
INV_X32 U_g18928 ( .A(g15606), .ZN(g18928) );
INV_X32 U_g18929 ( .A(g15609), .ZN(g18929) );
INV_X32 U_g18930 ( .A(g15612), .ZN(g18930) );
INV_X32 U_g18931 ( .A(g15615), .ZN(g18931) );
INV_X32 U_I24966 ( .A(g14863), .ZN(I24966) );
INV_X32 U_g18932 ( .A(I24966), .ZN(g18932) );
INV_X32 U_g18933 ( .A(g15625), .ZN(g18933) );
INV_X32 U_g18934 ( .A(g15628), .ZN(g18934) );
INV_X32 U_g18935 ( .A(g15631), .ZN(g18935) );
INV_X32 U_g18936 ( .A(g15635), .ZN(g18936) );
INV_X32 U_I24973 ( .A(g15003), .ZN(I24973) );
INV_X32 U_g18937 ( .A(I24973), .ZN(g18937) );
INV_X32 U_g18938 ( .A(g15641), .ZN(g18938) );
INV_X32 U_g18939 ( .A(g15644), .ZN(g18939) );
INV_X32 U_g18940 ( .A(g15647), .ZN(g18940) );
INV_X32 U_g18941 ( .A(g15652), .ZN(g18941) );
INV_X32 U_g18943 ( .A(g15655), .ZN(g18943) );
INV_X32 U_I24982 ( .A(g14347), .ZN(I24982) );
INV_X32 U_g18944 ( .A(I24982), .ZN(g18944) );
INV_X32 U_g18945 ( .A(g15667), .ZN(g18945) );
INV_X32 U_g18946 ( .A(g15672), .ZN(g18946) );
INV_X32 U_g18947 ( .A(g15675), .ZN(g18947) );
INV_X32 U_g18948 ( .A(g15682), .ZN(g18948) );
INV_X32 U_g18949 ( .A(g15685), .ZN(g18949) );
INV_X32 U_g18950 ( .A(g15688), .ZN(g18950) );
INV_X32 U_g18951 ( .A(g15691), .ZN(g18951) );
INV_X32 U_I24992 ( .A(g14936), .ZN(I24992) );
INV_X32 U_g18952 ( .A(I24992), .ZN(g18952) );
INV_X32 U_g18953 ( .A(g15701), .ZN(g18953) );
INV_X32 U_g18954 ( .A(g15704), .ZN(g18954) );
INV_X32 U_g18955 ( .A(g15707), .ZN(g18955) );
INV_X32 U_g18956 ( .A(g15711), .ZN(g18956) );
INV_X32 U_g18958 ( .A(g15714), .ZN(g18958) );
INV_X32 U_I25001 ( .A(g14244), .ZN(I25001) );
INV_X32 U_g18959 ( .A(I25001), .ZN(g18959) );
INV_X32 U_I25004 ( .A(g14459), .ZN(I25004) );
INV_X32 U_g18960 ( .A(I25004), .ZN(g18960) );
INV_X32 U_g18961 ( .A(g15726), .ZN(g18961) );
INV_X32 U_g18962 ( .A(g15731), .ZN(g18962) );
INV_X32 U_g18963 ( .A(g15734), .ZN(g18963) );
INV_X32 U_g18964 ( .A(g15741), .ZN(g18964) );
INV_X32 U_g18965 ( .A(g15744), .ZN(g18965) );
INV_X32 U_g18966 ( .A(g15747), .ZN(g18966) );
INV_X32 U_g18967 ( .A(g15750), .ZN(g18967) );
INV_X32 U_I25015 ( .A(g14158), .ZN(I25015) );
INV_X32 U_g18969 ( .A(I25015), .ZN(g18969) );
INV_X32 U_I25018 ( .A(g14366), .ZN(I25018) );
INV_X32 U_g18970 ( .A(I25018), .ZN(g18970) );
INV_X32 U_I25021 ( .A(g14546), .ZN(I25021) );
INV_X32 U_g18971 ( .A(I25021), .ZN(g18971) );
INV_X32 U_g18972 ( .A(g15766), .ZN(g18972) );
INV_X32 U_g18973 ( .A(g15771), .ZN(g18973) );
INV_X32 U_g18974 ( .A(g15774), .ZN(g18974) );
INV_X32 U_g18976 ( .A(g15777), .ZN(g18976) );
INV_X32 U_I25037 ( .A(g14071), .ZN(I25037) );
INV_X32 U_g18981 ( .A(I25037), .ZN(g18981) );
INV_X32 U_I25041 ( .A(g14895), .ZN(I25041) );
INV_X32 U_g18983 ( .A(I25041), .ZN(g18983) );
INV_X32 U_I25044 ( .A(g14273), .ZN(I25044) );
INV_X32 U_g18984 ( .A(I25044), .ZN(g18984) );
INV_X32 U_I25047 ( .A(g14478), .ZN(I25047) );
INV_X32 U_g18985 ( .A(I25047), .ZN(g18985) );
INV_X32 U_I25050 ( .A(g14601), .ZN(I25050) );
INV_X32 U_g18986 ( .A(I25050), .ZN(g18986) );
INV_X32 U_g18987 ( .A(g15794), .ZN(g18987) );
INV_X32 U_I25054 ( .A(g14837), .ZN(I25054) );
INV_X32 U_g18988 ( .A(I25054), .ZN(g18988) );
INV_X32 U_I25057 ( .A(g14186), .ZN(I25057) );
INV_X32 U_g18989 ( .A(I25057), .ZN(g18989) );
INV_X32 U_I25061 ( .A(g14976), .ZN(I25061) );
INV_X32 U_g18991 ( .A(I25061), .ZN(g18991) );
INV_X32 U_I25064 ( .A(g14395), .ZN(I25064) );
INV_X32 U_g18992 ( .A(I25064), .ZN(g18992) );
INV_X32 U_I25067 ( .A(g14565), .ZN(I25067) );
INV_X32 U_g18993 ( .A(I25067), .ZN(g18993) );
INV_X32 U_I25071 ( .A(g14910), .ZN(I25071) );
INV_X32 U_g18995 ( .A(I25071), .ZN(g18995) );
INV_X32 U_I25074 ( .A(g14301), .ZN(I25074) );
INV_X32 U_g18996 ( .A(I25074), .ZN(g18996) );
INV_X32 U_I25078 ( .A(g15065), .ZN(I25078) );
INV_X32 U_g18998 ( .A(I25078), .ZN(g18998) );
INV_X32 U_I25081 ( .A(g14507), .ZN(I25081) );
INV_X32 U_g18999 ( .A(I25081), .ZN(g18999) );
INV_X32 U_I25084 ( .A(g14885), .ZN(I25084) );
INV_X32 U_g19000 ( .A(I25084), .ZN(g19000) );
INV_X32 U_g19001 ( .A(g14071), .ZN(g19001) );
INV_X32 U_I25089 ( .A(g14991), .ZN(I25089) );
INV_X32 U_g19008 ( .A(I25089), .ZN(g19008) );
INV_X32 U_I25092 ( .A(g14423), .ZN(I25092) );
INV_X32 U_g19009 ( .A(I25092), .ZN(g19009) );
INV_X32 U_I25096 ( .A(g15161), .ZN(I25096) );
INV_X32 U_g19011 ( .A(I25096), .ZN(g19011) );
INV_X32 U_I25099 ( .A(g19000), .ZN(I25099) );
INV_X32 U_g19012 ( .A(I25099), .ZN(g19012) );
INV_X32 U_I25102 ( .A(g18944), .ZN(I25102) );
INV_X32 U_g19013 ( .A(I25102), .ZN(g19013) );
INV_X32 U_I25105 ( .A(g18959), .ZN(I25105) );
INV_X32 U_g19014 ( .A(I25105), .ZN(g19014) );
INV_X32 U_I25108 ( .A(g18969), .ZN(I25108) );
INV_X32 U_g19015 ( .A(I25108), .ZN(g19015) );
INV_X32 U_I25111 ( .A(g18981), .ZN(I25111) );
INV_X32 U_g19016 ( .A(I25111), .ZN(g19016) );
INV_X32 U_I25114 ( .A(g18983), .ZN(I25114) );
INV_X32 U_g19017 ( .A(I25114), .ZN(g19017) );
INV_X32 U_I25117 ( .A(g18988), .ZN(I25117) );
INV_X32 U_g19018 ( .A(I25117), .ZN(g19018) );
INV_X32 U_I25120 ( .A(g18869), .ZN(I25120) );
INV_X32 U_g19019 ( .A(I25120), .ZN(g19019) );
INV_X32 U_I25123 ( .A(g18890), .ZN(I25123) );
INV_X32 U_g19020 ( .A(I25123), .ZN(g19020) );
INV_X32 U_I25126 ( .A(g16858), .ZN(I25126) );
INV_X32 U_g19021 ( .A(I25126), .ZN(g19021) );
INV_X32 U_I25129 ( .A(g16813), .ZN(I25129) );
INV_X32 U_g19022 ( .A(I25129), .ZN(g19022) );
INV_X32 U_I25132 ( .A(g16862), .ZN(I25132) );
INV_X32 U_g19023 ( .A(I25132), .ZN(g19023) );
INV_X32 U_I25135 ( .A(g16506), .ZN(I25135) );
INV_X32 U_g19024 ( .A(I25135), .ZN(g19024) );
INV_X32 U_I25138 ( .A(g18960), .ZN(I25138) );
INV_X32 U_g19025 ( .A(I25138), .ZN(g19025) );
INV_X32 U_I25141 ( .A(g18970), .ZN(I25141) );
INV_X32 U_g19026 ( .A(I25141), .ZN(g19026) );
INV_X32 U_I25144 ( .A(g18984), .ZN(I25144) );
INV_X32 U_g19027 ( .A(I25144), .ZN(g19027) );
INV_X32 U_I25147 ( .A(g18989), .ZN(I25147) );
INV_X32 U_g19028 ( .A(I25147), .ZN(g19028) );
INV_X32 U_I25150 ( .A(g18991), .ZN(I25150) );
INV_X32 U_g19029 ( .A(I25150), .ZN(g19029) );
INV_X32 U_I25153 ( .A(g18995), .ZN(I25153) );
INV_X32 U_g19030 ( .A(I25153), .ZN(g19030) );
INV_X32 U_I25156 ( .A(g18895), .ZN(I25156) );
INV_X32 U_g19031 ( .A(I25156), .ZN(g19031) );
INV_X32 U_I25159 ( .A(g18913), .ZN(I25159) );
INV_X32 U_g19032 ( .A(I25159), .ZN(g19032) );
INV_X32 U_I25162 ( .A(g16863), .ZN(I25162) );
INV_X32 U_g19033 ( .A(I25162), .ZN(g19033) );
INV_X32 U_I25165 ( .A(g16831), .ZN(I25165) );
INV_X32 U_g19034 ( .A(I25165), .ZN(g19034) );
INV_X32 U_I25168 ( .A(g16877), .ZN(I25168) );
INV_X32 U_g19035 ( .A(I25168), .ZN(g19035) );
INV_X32 U_I25171 ( .A(g16528), .ZN(I25171) );
INV_X32 U_g19036 ( .A(I25171), .ZN(g19036) );
INV_X32 U_I25174 ( .A(g18971), .ZN(I25174) );
INV_X32 U_g19037 ( .A(I25174), .ZN(g19037) );
INV_X32 U_I25177 ( .A(g18985), .ZN(I25177) );
INV_X32 U_g19038 ( .A(I25177), .ZN(g19038) );
INV_X32 U_I25180 ( .A(g18992), .ZN(I25180) );
INV_X32 U_g19039 ( .A(I25180), .ZN(g19039) );
INV_X32 U_I25183 ( .A(g18996), .ZN(I25183) );
INV_X32 U_g19040 ( .A(I25183), .ZN(g19040) );
INV_X32 U_I25186 ( .A(g18998), .ZN(I25186) );
INV_X32 U_g19041 ( .A(I25186), .ZN(g19041) );
INV_X32 U_I25189 ( .A(g19008), .ZN(I25189) );
INV_X32 U_g19042 ( .A(I25189), .ZN(g19042) );
INV_X32 U_I25192 ( .A(g18918), .ZN(I25192) );
INV_X32 U_g19043 ( .A(I25192), .ZN(g19043) );
INV_X32 U_I25195 ( .A(g18932), .ZN(I25195) );
INV_X32 U_g19044 ( .A(I25195), .ZN(g19044) );
INV_X32 U_I25198 ( .A(g16878), .ZN(I25198) );
INV_X32 U_g19045 ( .A(I25198), .ZN(g19045) );
INV_X32 U_I25201 ( .A(g16843), .ZN(I25201) );
INV_X32 U_g19046 ( .A(I25201), .ZN(g19046) );
INV_X32 U_I25204 ( .A(g16905), .ZN(I25204) );
INV_X32 U_g19047 ( .A(I25204), .ZN(g19047) );
INV_X32 U_I25207 ( .A(g16559), .ZN(I25207) );
INV_X32 U_g19048 ( .A(I25207), .ZN(g19048) );
INV_X32 U_I25210 ( .A(g18986), .ZN(I25210) );
INV_X32 U_g19049 ( .A(I25210), .ZN(g19049) );
INV_X32 U_I25213 ( .A(g18993), .ZN(I25213) );
INV_X32 U_g19050 ( .A(I25213), .ZN(g19050) );
INV_X32 U_I25216 ( .A(g18999), .ZN(I25216) );
INV_X32 U_g19051 ( .A(I25216), .ZN(g19051) );
INV_X32 U_I25219 ( .A(g19009), .ZN(I25219) );
INV_X32 U_g19052 ( .A(I25219), .ZN(g19052) );
INV_X32 U_I25222 ( .A(g19011), .ZN(I25222) );
INV_X32 U_g19053 ( .A(I25222), .ZN(g19053) );
INV_X32 U_I25225 ( .A(g16514), .ZN(I25225) );
INV_X32 U_g19054 ( .A(I25225), .ZN(g19054) );
INV_X32 U_I25228 ( .A(g18937), .ZN(I25228) );
INV_X32 U_g19055 ( .A(I25228), .ZN(g19055) );
INV_X32 U_I25231 ( .A(g18952), .ZN(I25231) );
INV_X32 U_g19056 ( .A(I25231), .ZN(g19056) );
INV_X32 U_I25234 ( .A(g16906), .ZN(I25234) );
INV_X32 U_g19057 ( .A(I25234), .ZN(g19057) );
INV_X32 U_I25237 ( .A(g16849), .ZN(I25237) );
INV_X32 U_g19058 ( .A(I25237), .ZN(g19058) );
INV_X32 U_I25240 ( .A(g16934), .ZN(I25240) );
INV_X32 U_g19059 ( .A(I25240), .ZN(g19059) );
INV_X32 U_I25243 ( .A(g17227), .ZN(I25243) );
INV_X32 U_g19060 ( .A(I25243), .ZN(g19060) );
INV_X32 U_I25246 ( .A(g17233), .ZN(I25246) );
INV_X32 U_g19061 ( .A(I25246), .ZN(g19061) );
INV_X32 U_I25249 ( .A(g17300), .ZN(I25249) );
INV_X32 U_g19062 ( .A(I25249), .ZN(g19062) );
INV_X32 U_I25253 ( .A(g17124), .ZN(I25253) );
INV_X32 U_g19064 ( .A(I25253), .ZN(g19064) );
INV_X32 U_g19070 ( .A(g18583), .ZN(g19070) );
INV_X32 U_I25258 ( .A(g16974), .ZN(I25258) );
INV_X32 U_g19075 ( .A(I25258), .ZN(g19075) );
INV_X32 U_g19078 ( .A(g18619), .ZN(g19078) );
INV_X32 U_I25264 ( .A(g17151), .ZN(I25264) );
INV_X32 U_g19081 ( .A(I25264), .ZN(g19081) );
INV_X32 U_I25272 ( .A(g17051), .ZN(I25272) );
INV_X32 U_g19091 ( .A(I25272), .ZN(g19091) );
INV_X32 U_g19096 ( .A(g18980), .ZN(g19096) );
INV_X32 U_I25283 ( .A(g17086), .ZN(I25283) );
INV_X32 U_g19098 ( .A(I25283), .ZN(g19098) );
INV_X32 U_I25294 ( .A(g17124), .ZN(I25294) );
INV_X32 U_g19105 ( .A(I25294), .ZN(g19105) );
INV_X32 U_I25303 ( .A(g17151), .ZN(I25303) );
INV_X32 U_g19110 ( .A(I25303), .ZN(g19110) );
INV_X32 U_I25308 ( .A(g16867), .ZN(I25308) );
INV_X32 U_g19113 ( .A(I25308), .ZN(g19113) );
INV_X32 U_I25315 ( .A(g16895), .ZN(I25315) );
INV_X32 U_g19118 ( .A(I25315), .ZN(g19118) );
INV_X32 U_I25320 ( .A(g16924), .ZN(I25320) );
INV_X32 U_g19125 ( .A(I25320), .ZN(g19125) );
INV_X32 U_I25325 ( .A(g16954), .ZN(I25325) );
INV_X32 U_g19132 ( .A(I25325), .ZN(g19132) );
INV_X32 U_I25334 ( .A(g17645), .ZN(I25334) );
INV_X32 U_g19145 ( .A(I25334), .ZN(g19145) );
INV_X32 U_I25338 ( .A(g17746), .ZN(I25338) );
INV_X32 U_g19147 ( .A(I25338), .ZN(g19147) );
INV_X32 U_I25344 ( .A(g17847), .ZN(I25344) );
INV_X32 U_g19151 ( .A(I25344), .ZN(g19151) );
INV_X32 U_I25351 ( .A(g17959), .ZN(I25351) );
INV_X32 U_g19156 ( .A(I25351), .ZN(g19156) );
INV_X32 U_I25355 ( .A(g18669), .ZN(I25355) );
INV_X32 U_g19158 ( .A(I25355), .ZN(g19158) );
INV_X32 U_I25358 ( .A(g18678), .ZN(I25358) );
INV_X32 U_g19159 ( .A(I25358), .ZN(g19159) );
INV_X32 U_I25365 ( .A(g18707), .ZN(I25365) );
INV_X32 U_g19164 ( .A(I25365), .ZN(g19164) );
INV_X32 U_I25371 ( .A(g18719), .ZN(I25371) );
INV_X32 U_g19168 ( .A(I25371), .ZN(g19168) );
INV_X32 U_I25374 ( .A(g18726), .ZN(I25374) );
INV_X32 U_g19169 ( .A(I25374), .ZN(g19169) );
INV_X32 U_I25377 ( .A(g18743), .ZN(I25377) );
INV_X32 U_g19170 ( .A(I25377), .ZN(g19170) );
INV_X32 U_I25383 ( .A(g18755), .ZN(I25383) );
INV_X32 U_g19174 ( .A(I25383), .ZN(g19174) );
INV_X32 U_I25386 ( .A(g18763), .ZN(I25386) );
INV_X32 U_g19175 ( .A(I25386), .ZN(g19175) );
INV_X32 U_I25389 ( .A(g18780), .ZN(I25389) );
INV_X32 U_g19176 ( .A(I25389), .ZN(g19176) );
INV_X32 U_I25395 ( .A(g18782), .ZN(I25395) );
INV_X32 U_g19180 ( .A(I25395), .ZN(g19180) );
INV_X32 U_I25399 ( .A(g18794), .ZN(I25399) );
INV_X32 U_g19182 ( .A(I25399), .ZN(g19182) );
INV_X32 U_I25402 ( .A(g18821), .ZN(I25402) );
INV_X32 U_g19183 ( .A(I25402), .ZN(g19183) );
INV_X32 U_I25406 ( .A(g18804), .ZN(I25406) );
INV_X32 U_g19185 ( .A(I25406), .ZN(g19185) );
INV_X32 U_I25412 ( .A(g18820), .ZN(I25412) );
INV_X32 U_g19189 ( .A(I25412), .ZN(g19189) );
INV_X32 U_I25415 ( .A(g18835), .ZN(I25415) );
INV_X32 U_g19190 ( .A(I25415), .ZN(g19190) );
INV_X32 U_I25423 ( .A(g18852), .ZN(I25423) );
INV_X32 U_g19196 ( .A(I25423), .ZN(g19196) );
INV_X32 U_I25426 ( .A(g18836), .ZN(I25426) );
INV_X32 U_g19197 ( .A(I25426), .ZN(g19197) );
INV_X32 U_I25429 ( .A(g18975), .ZN(I25429) );
INV_X32 U_g19198 ( .A(I25429), .ZN(g19198) );
INV_X32 U_I25432 ( .A(g18837), .ZN(I25432) );
INV_X32 U_g19199 ( .A(I25432), .ZN(g19199) );
INV_X32 U_I25442 ( .A(g18866), .ZN(I25442) );
INV_X32 U_g19207 ( .A(I25442), .ZN(g19207) );
INV_X32 U_I25445 ( .A(g18968), .ZN(I25445) );
INV_X32 U_g19208 ( .A(I25445), .ZN(g19208) );
INV_X32 U_I25456 ( .A(g18883), .ZN(I25456) );
INV_X32 U_g19217 ( .A(I25456), .ZN(g19217) );
INV_X32 U_I25459 ( .A(g18867), .ZN(I25459) );
INV_X32 U_g19218 ( .A(I25459), .ZN(g19218) );
INV_X32 U_I25463 ( .A(g18868), .ZN(I25463) );
INV_X32 U_g19220 ( .A(I25463), .ZN(g19220) );
INV_X32 U_I25474 ( .A(g18885), .ZN(I25474) );
INV_X32 U_g19229 ( .A(I25474), .ZN(g19229) );
INV_X32 U_I25486 ( .A(g18754), .ZN(I25486) );
INV_X32 U_g19237 ( .A(I25486), .ZN(g19237) );
INV_X32 U_I25489 ( .A(g18906), .ZN(I25489) );
INV_X32 U_g19238 ( .A(I25489), .ZN(g19238) );
INV_X32 U_I25492 ( .A(g18907), .ZN(I25492) );
INV_X32 U_g19239 ( .A(I25492), .ZN(g19239) );
INV_X32 U_I25506 ( .A(g18781), .ZN(I25506) );
INV_X32 U_g19247 ( .A(I25506), .ZN(g19247) );
INV_X32 U_I25510 ( .A(g18542), .ZN(I25510) );
INV_X32 U_g19249 ( .A(I25510), .ZN(g19249) );
INV_X32 U_g19251 ( .A(g16540), .ZN(g19251) );
INV_X32 U_I25525 ( .A(g18803), .ZN(I25525) );
INV_X32 U_g19258 ( .A(I25525), .ZN(g19258) );
INV_X32 U_I25528 ( .A(g18942), .ZN(I25528) );
INV_X32 U_g19259 ( .A(I25528), .ZN(g19259) );
INV_X32 U_g19265 ( .A(g16572), .ZN(g19265) );
INV_X32 U_I25557 ( .A(g18957), .ZN(I25557) );
INV_X32 U_g19270 ( .A(I25557), .ZN(g19270) );
INV_X32 U_I25567 ( .A(g17186), .ZN(I25567) );
INV_X32 U_g19272 ( .A(I25567), .ZN(g19272) );
INV_X32 U_g19280 ( .A(g16596), .ZN(g19280) );
INV_X32 U_g19287 ( .A(g16608), .ZN(g19287) );
INV_X32 U_I25612 ( .A(g17197), .ZN(I25612) );
INV_X32 U_g19291 ( .A(I25612), .ZN(g19291) );
INV_X32 U_g19299 ( .A(g16616), .ZN(g19299) );
INV_X32 U_g19301 ( .A(g16622), .ZN(g19301) );
INV_X32 U_g19302 ( .A(g17025), .ZN(g19302) );
INV_X32 U_g19305 ( .A(g16626), .ZN(g19305) );
INV_X32 U_I25660 ( .A(g17204), .ZN(I25660) );
INV_X32 U_g19309 ( .A(I25660), .ZN(g19309) );
INV_X32 U_g19319 ( .A(g16633), .ZN(g19319) );
INV_X32 U_g19322 ( .A(g16636), .ZN(g19322) );
INV_X32 U_g19323 ( .A(g17059), .ZN(g19323) );
INV_X32 U_g19326 ( .A(g16640), .ZN(g19326) );
INV_X32 U_I25717 ( .A(g17209), .ZN(I25717) );
INV_X32 U_g19330 ( .A(I25717), .ZN(g19330) );
INV_X32 U_I25728 ( .A(g17118), .ZN(I25728) );
INV_X32 U_g19335 ( .A(I25728), .ZN(g19335) );
INV_X32 U_g19346 ( .A(g16644), .ZN(g19346) );
INV_X32 U_g19349 ( .A(g16647), .ZN(g19349) );
INV_X32 U_g19350 ( .A(g17094), .ZN(g19350) );
INV_X32 U_g19353 ( .A(g16651), .ZN(g19353) );
INV_X32 U_I25768 ( .A(g17139), .ZN(I25768) );
INV_X32 U_g19358 ( .A(I25768), .ZN(g19358) );
INV_X32 U_I25778 ( .A(g17145), .ZN(I25778) );
INV_X32 U_g19369 ( .A(I25778), .ZN(g19369) );
INV_X32 U_g19380 ( .A(g16656), .ZN(g19380) );
INV_X32 U_g19383 ( .A(g16659), .ZN(g19383) );
INV_X32 U_g19384 ( .A(g17132), .ZN(g19384) );
INV_X32 U_g19387 ( .A(g16567), .ZN(g19387) );
INV_X32 U_g19388 ( .A(g17139), .ZN(g19388) );
INV_X32 U_I25816 ( .A(g17162), .ZN(I25816) );
INV_X32 U_g19390 ( .A(I25816), .ZN(g19390) );
INV_X32 U_I25826 ( .A(g17168), .ZN(I25826) );
INV_X32 U_g19401 ( .A(I25826), .ZN(g19401) );
INV_X32 U_g19412 ( .A(g16673), .ZN(g19412) );
INV_X32 U_g19415 ( .A(g16676), .ZN(g19415) );
INV_X32 U_g19417 ( .A(g16591), .ZN(g19417) );
INV_X32 U_g19418 ( .A(g17162), .ZN(g19418) );
INV_X32 U_I25862 ( .A(g17177), .ZN(I25862) );
INV_X32 U_g19420 ( .A(I25862), .ZN(g19420) );
INV_X32 U_I25872 ( .A(g17183), .ZN(I25872) );
INV_X32 U_g19431 ( .A(I25872), .ZN(g19431) );
INV_X32 U_g19441 ( .A(g17213), .ZN(g19441) );
INV_X32 U_g19444 ( .A(g17985), .ZN(g19444) );
INV_X32 U_g19448 ( .A(g16694), .ZN(g19448) );
INV_X32 U_g19452 ( .A(g16702), .ZN(g19452) );
INV_X32 U_g19454 ( .A(g16611), .ZN(g19454) );
INV_X32 U_g19455 ( .A(g17177), .ZN(g19455) );
INV_X32 U_I25904 ( .A(g17194), .ZN(I25904) );
INV_X32 U_g19457 ( .A(I25904), .ZN(g19457) );
INV_X32 U_g19467 ( .A(g16719), .ZN(g19467) );
INV_X32 U_g19468 ( .A(g17216), .ZN(g19468) );
INV_X32 U_g19471 ( .A(g18102), .ZN(g19471) );
INV_X32 U_g19475 ( .A(g16725), .ZN(g19475) );
INV_X32 U_g19479 ( .A(g16733), .ZN(g19479) );
INV_X32 U_g19481 ( .A(g16629), .ZN(g19481) );
INV_X32 U_g19482 ( .A(g17194), .ZN(g19482) );
INV_X32 U_g19483 ( .A(g16758), .ZN(g19483) );
INV_X32 U_g19484 ( .A(g16867), .ZN(g19484) );
INV_X32 U_g19490 ( .A(g16761), .ZN(g19490) );
INV_X32 U_g19491 ( .A(g17219), .ZN(g19491) );
INV_X32 U_g19494 ( .A(g18218), .ZN(g19494) );
INV_X32 U_g19498 ( .A(g16767), .ZN(g19498) );
INV_X32 U_g19502 ( .A(g16775), .ZN(g19502) );
INV_X32 U_g19504 ( .A(g16785), .ZN(g19504) );
INV_X32 U_g19505 ( .A(g16895), .ZN(g19505) );
INV_X32 U_g19511 ( .A(g16788), .ZN(g19511) );
INV_X32 U_g19512 ( .A(g17221), .ZN(g19512) );
INV_X32 U_g19515 ( .A(g18325), .ZN(g19515) );
INV_X32 U_g19519 ( .A(g16794), .ZN(g19519) );
INV_X32 U_g19523 ( .A(g16814), .ZN(g19523) );
INV_X32 U_g19524 ( .A(g16924), .ZN(g19524) );
INV_X32 U_g19530 ( .A(g16817), .ZN(g19530) );
INV_X32 U_g19533 ( .A(g16832), .ZN(g19533) );
INV_X32 U_g19534 ( .A(g16954), .ZN(g19534) );
INV_X32 U_I25966 ( .A(g16654), .ZN(I25966) );
INV_X32 U_g19543 ( .A(I25966), .ZN(g19543) );
INV_X32 U_I25971 ( .A(g16671), .ZN(I25971) );
INV_X32 U_g19546 ( .A(I25971), .ZN(g19546) );
INV_X32 U_I25977 ( .A(g16692), .ZN(I25977) );
INV_X32 U_g19550 ( .A(I25977), .ZN(g19550) );
INV_X32 U_I25985 ( .A(g16718), .ZN(I25985) );
INV_X32 U_g19556 ( .A(I25985), .ZN(g19556) );
INV_X32 U_I25994 ( .A(g16860), .ZN(I25994) );
INV_X32 U_g19563 ( .A(I25994), .ZN(g19563) );
INV_X32 U_I26006 ( .A(g16866), .ZN(I26006) );
INV_X32 U_g19573 ( .A(I26006), .ZN(g19573) );
INV_X32 U_g19577 ( .A(g16881), .ZN(g19577) );
INV_X32 U_g19578 ( .A(g16884), .ZN(g19578) );
INV_X32 U_I26025 ( .A(g16803), .ZN(I26025) );
INV_X32 U_g19595 ( .A(I26025), .ZN(g19595) );
INV_X32 U_I26028 ( .A(g16566), .ZN(I26028) );
INV_X32 U_g19596 ( .A(I26028), .ZN(g19596) );
INV_X32 U_g19607 ( .A(g16910), .ZN(g19607) );
INV_X32 U_g19608 ( .A(g16913), .ZN(g19608) );
INV_X32 U_I26051 ( .A(g16824), .ZN(I26051) );
INV_X32 U_g19622 ( .A(I26051), .ZN(g19622) );
INV_X32 U_g19640 ( .A(g16940), .ZN(g19640) );
INV_X32 U_g19641 ( .A(g16943), .ZN(g19641) );
INV_X32 U_I26078 ( .A(g16835), .ZN(I26078) );
INV_X32 U_g19652 ( .A(I26078), .ZN(g19652) );
INV_X32 U_I26085 ( .A(g18085), .ZN(I26085) );
INV_X32 U_g19657 ( .A(I26085), .ZN(g19657) );
INV_X32 U_g19680 ( .A(g16971), .ZN(g19680) );
INV_X32 U_g19681 ( .A(g16974), .ZN(g19681) );
INV_X32 U_I26112 ( .A(g16844), .ZN(I26112) );
INV_X32 U_g19689 ( .A(I26112), .ZN(g19689) );
INV_X32 U_I26115 ( .A(g16845), .ZN(I26115) );
INV_X32 U_g19690 ( .A(I26115), .ZN(g19690) );
INV_X32 U_I26123 ( .A(g17503), .ZN(I26123) );
INV_X32 U_g19696 ( .A(I26123), .ZN(g19696) );
INV_X32 U_I26134 ( .A(g18201), .ZN(I26134) );
INV_X32 U_g19705 ( .A(I26134), .ZN(g19705) );
INV_X32 U_I26154 ( .A(g16851), .ZN(I26154) );
INV_X32 U_g19725 ( .A(I26154), .ZN(g19725) );
INV_X32 U_I26171 ( .A(g17594), .ZN(I26171) );
INV_X32 U_g19740 ( .A(I26171), .ZN(g19740) );
INV_X32 U_I26182 ( .A(g18308), .ZN(I26182) );
INV_X32 U_g19749 ( .A(I26182), .ZN(g19749) );
INV_X32 U_I26195 ( .A(g16853), .ZN(I26195) );
INV_X32 U_g19762 ( .A(I26195), .ZN(g19762) );
INV_X32 U_I26198 ( .A(g16854), .ZN(I26198) );
INV_X32 U_g19763 ( .A(I26198), .ZN(g19763) );
INV_X32 U_I26220 ( .A(g17691), .ZN(I26220) );
INV_X32 U_g19783 ( .A(I26220), .ZN(g19783) );
INV_X32 U_I26231 ( .A(g18401), .ZN(I26231) );
INV_X32 U_g19792 ( .A(I26231), .ZN(g19792) );
INV_X32 U_I26237 ( .A(g16857), .ZN(I26237) );
INV_X32 U_g19798 ( .A(I26237), .ZN(g19798) );
INV_X32 U_I26266 ( .A(g17791), .ZN(I26266) );
INV_X32 U_g19825 ( .A(I26266), .ZN(g19825) );
INV_X32 U_g19830 ( .A(g18886), .ZN(g19830) );
INV_X32 U_I26276 ( .A(g16861), .ZN(I26276) );
INV_X32 U_g19838 ( .A(I26276), .ZN(g19838) );
INV_X32 U_I26334 ( .A(g18977), .ZN(I26334) );
INV_X32 U_g19890 ( .A(I26334), .ZN(g19890) );
INV_X32 U_I26337 ( .A(g16880), .ZN(I26337) );
INV_X32 U_g19893 ( .A(I26337), .ZN(g19893) );
INV_X32 U_I26340 ( .A(g17025), .ZN(I26340) );
INV_X32 U_g19894 ( .A(I26340), .ZN(g19894) );
INV_X32 U_I26365 ( .A(g18626), .ZN(I26365) );
INV_X32 U_g19915 ( .A(I26365), .ZN(g19915) );
INV_X32 U_g19918 ( .A(g18646), .ZN(g19918) );
INV_X32 U_I26369 ( .A(g17059), .ZN(I26369) );
INV_X32 U_g19919 ( .A(I26369), .ZN(g19919) );
INV_X32 U_g19933 ( .A(g18548), .ZN(g19933) );
INV_X32 U_I26388 ( .A(g17094), .ZN(I26388) );
INV_X32 U_g19934 ( .A(I26388), .ZN(g19934) );
INV_X32 U_I26401 ( .A(g17012), .ZN(I26401) );
INV_X32 U_g19945 ( .A(I26401), .ZN(g19945) );
INV_X32 U_g19948 ( .A(g17896), .ZN(g19948) );
INV_X32 U_g19950 ( .A(g18598), .ZN(g19950) );
INV_X32 U_I26407 ( .A(g17132), .ZN(I26407) );
INV_X32 U_g19951 ( .A(I26407), .ZN(g19951) );
INV_X32 U_I26413 ( .A(g16643), .ZN(I26413) );
INV_X32 U_g19957 ( .A(I26413), .ZN(g19957) );
INV_X32 U_I26420 ( .A(g17042), .ZN(I26420) );
INV_X32 U_g19972 ( .A(I26420), .ZN(g19972) );
INV_X32 U_g19975 ( .A(g18007), .ZN(g19975) );
INV_X32 U_g19977 ( .A(g18630), .ZN(g19977) );
INV_X32 U_I26426 ( .A(g16536), .ZN(I26426) );
INV_X32 U_g19978 ( .A(I26426), .ZN(g19978) );
INV_X32 U_I26437 ( .A(g16655), .ZN(I26437) );
INV_X32 U_g19987 ( .A(I26437), .ZN(g19987) );
INV_X32 U_I26444 ( .A(g17076), .ZN(I26444) );
INV_X32 U_g20002 ( .A(I26444), .ZN(g20002) );
INV_X32 U_g20005 ( .A(g18124), .ZN(g20005) );
INV_X32 U_g20007 ( .A(g18639), .ZN(g20007) );
INV_X32 U_I26458 ( .A(g17985), .ZN(I26458) );
INV_X32 U_g20016 ( .A(I26458), .ZN(g20016) );
INV_X32 U_I26469 ( .A(g16672), .ZN(I26469) );
INV_X32 U_g20025 ( .A(I26469), .ZN(g20025) );
INV_X32 U_I26476 ( .A(g17111), .ZN(I26476) );
INV_X32 U_g20040 ( .A(I26476), .ZN(g20040) );
INV_X32 U_g20043 ( .A(g18240), .ZN(g20043) );
INV_X32 U_I26481 ( .A(g18590), .ZN(I26481) );
INV_X32 U_g20045 ( .A(I26481), .ZN(g20045) );
INV_X32 U_I26494 ( .A(g18102), .ZN(I26494) );
INV_X32 U_g20058 ( .A(I26494), .ZN(g20058) );
INV_X32 U_I26505 ( .A(g16693), .ZN(I26505) );
INV_X32 U_g20067 ( .A(I26505), .ZN(g20067) );
INV_X32 U_I26512 ( .A(g16802), .ZN(I26512) );
INV_X32 U_g20082 ( .A(I26512), .ZN(g20082) );
INV_X32 U_g20083 ( .A(g17968), .ZN(g20083) );
INV_X32 U_I26535 ( .A(g18218), .ZN(I26535) );
INV_X32 U_g20099 ( .A(I26535), .ZN(g20099) );
INV_X32 U_I26545 ( .A(g16823), .ZN(I26545) );
INV_X32 U_g20105 ( .A(I26545), .ZN(g20105) );
INV_X32 U_I26574 ( .A(g18325), .ZN(I26574) );
INV_X32 U_g20124 ( .A(I26574), .ZN(g20124) );
INV_X32 U_g20127 ( .A(g18623), .ZN(g20127) );
INV_X32 U_g20140 ( .A(g16830), .ZN(g20140) );
INV_X32 U_g20163 ( .A(g17973), .ZN(g20163) );
INV_X32 U_I26612 ( .A(g17645), .ZN(I26612) );
INV_X32 U_g20164 ( .A(I26612), .ZN(g20164) );
INV_X32 U_g20178 ( .A(g16842), .ZN(g20178) );
INV_X32 U_g20193 ( .A(g18691), .ZN(g20193) );
INV_X32 U_I26642 ( .A(g17746), .ZN(I26642) );
INV_X32 U_g20198 ( .A(I26642), .ZN(g20198) );
INV_X32 U_g20212 ( .A(g16848), .ZN(g20212) );
INV_X32 U_g20223 ( .A(g18727), .ZN(g20223) );
INV_X32 U_I26664 ( .A(g17847), .ZN(I26664) );
INV_X32 U_g20228 ( .A(I26664), .ZN(g20228) );
INV_X32 U_g20242 ( .A(g16852), .ZN(g20242) );
INV_X32 U_g20250 ( .A(g18764), .ZN(g20250) );
INV_X32 U_I26679 ( .A(g17959), .ZN(I26679) );
INV_X32 U_g20255 ( .A(I26679), .ZN(g20255) );
INV_X32 U_g20269 ( .A(g17230), .ZN(g20269) );
INV_X32 U_g20273 ( .A(g18795), .ZN(g20273) );
INV_X32 U_g20278 ( .A(g17237), .ZN(g20278) );
INV_X32 U_g20279 ( .A(g17240), .ZN(g20279) );
INV_X32 U_g20281 ( .A(g17243), .ZN(g20281) );
INV_X32 U_g20286 ( .A(g17249), .ZN(g20286) );
INV_X32 U_g20287 ( .A(g17252), .ZN(g20287) );
INV_X32 U_g20288 ( .A(g17255), .ZN(g20288) );
INV_X32 U_g20289 ( .A(g17259), .ZN(g20289) );
INV_X32 U_g20290 ( .A(g17262), .ZN(g20290) );
INV_X32 U_g20292 ( .A(g17265), .ZN(g20292) );
INV_X32 U_I26714 ( .A(g17720), .ZN(I26714) );
INV_X32 U_g20295 ( .A(I26714), .ZN(g20295) );
INV_X32 U_g20296 ( .A(g17272), .ZN(g20296) );
INV_X32 U_g20297 ( .A(g17275), .ZN(g20297) );
INV_X32 U_g20298 ( .A(g17278), .ZN(g20298) );
INV_X32 U_g20302 ( .A(g17282), .ZN(g20302) );
INV_X32 U_g20303 ( .A(g17285), .ZN(g20303) );
INV_X32 U_g20304 ( .A(g17288), .ZN(g20304) );
INV_X32 U_g20305 ( .A(g17291), .ZN(g20305) );
INV_X32 U_g20306 ( .A(g17294), .ZN(g20306) );
INV_X32 U_g20308 ( .A(g17297), .ZN(g20308) );
INV_X32 U_g20311 ( .A(g17304), .ZN(g20311) );
INV_X32 U_g20312 ( .A(g17307), .ZN(g20312) );
INV_X32 U_g20313 ( .A(g17310), .ZN(g20313) );
INV_X32 U_g20315 ( .A(g17315), .ZN(g20315) );
INV_X32 U_g20316 ( .A(g17318), .ZN(g20316) );
INV_X32 U_g20317 ( .A(g17321), .ZN(g20317) );
INV_X32 U_g20321 ( .A(g17324), .ZN(g20321) );
INV_X32 U_g20322 ( .A(g17327), .ZN(g20322) );
INV_X32 U_g20323 ( .A(g17330), .ZN(g20323) );
INV_X32 U_g20324 ( .A(g17333), .ZN(g20324) );
INV_X32 U_g20325 ( .A(g17336), .ZN(g20325) );
INV_X32 U_g20327 ( .A(g17342), .ZN(g20327) );
INV_X32 U_g20328 ( .A(g17345), .ZN(g20328) );
INV_X32 U_g20329 ( .A(g17348), .ZN(g20329) );
INV_X32 U_g20330 ( .A(g17354), .ZN(g20330) );
INV_X32 U_g20331 ( .A(g17357), .ZN(g20331) );
INV_X32 U_g20332 ( .A(g17360), .ZN(g20332) );
INV_X32 U_g20334 ( .A(g17363), .ZN(g20334) );
INV_X32 U_g20335 ( .A(g17366), .ZN(g20335) );
INV_X32 U_g20336 ( .A(g17369), .ZN(g20336) );
INV_X32 U_g20340 ( .A(g17372), .ZN(g20340) );
INV_X32 U_g20341 ( .A(g17375), .ZN(g20341) );
INV_X32 U_g20342 ( .A(g17378), .ZN(g20342) );
INV_X32 U_g20344 ( .A(g17384), .ZN(g20344) );
INV_X32 U_g20345 ( .A(g17387), .ZN(g20345) );
INV_X32 U_g20346 ( .A(g17390), .ZN(g20346) );
INV_X32 U_g20347 ( .A(g17399), .ZN(g20347) );
INV_X32 U_g20348 ( .A(g17402), .ZN(g20348) );
INV_X32 U_g20349 ( .A(g17405), .ZN(g20349) );
INV_X32 U_g20350 ( .A(g17410), .ZN(g20350) );
INV_X32 U_g20351 ( .A(g17413), .ZN(g20351) );
INV_X32 U_g20352 ( .A(g17416), .ZN(g20352) );
INV_X32 U_g20354 ( .A(g17419), .ZN(g20354) );
INV_X32 U_g20355 ( .A(g17422), .ZN(g20355) );
INV_X32 U_g20356 ( .A(g17425), .ZN(g20356) );
INV_X32 U_I26777 ( .A(g17222), .ZN(I26777) );
INV_X32 U_g20360 ( .A(I26777), .ZN(g20360) );
INV_X32 U_g20361 ( .A(g17430), .ZN(g20361) );
INV_X32 U_g20362 ( .A(g17433), .ZN(g20362) );
INV_X32 U_g20363 ( .A(g17436), .ZN(g20363) );
INV_X32 U_g20364 ( .A(g17439), .ZN(g20364) );
INV_X32 U_g20365 ( .A(g17442), .ZN(g20365) );
INV_X32 U_g20366 ( .A(g17451), .ZN(g20366) );
INV_X32 U_g20367 ( .A(g17454), .ZN(g20367) );
INV_X32 U_g20368 ( .A(g17457), .ZN(g20368) );
INV_X32 U_g20369 ( .A(g17465), .ZN(g20369) );
INV_X32 U_g20370 ( .A(g17468), .ZN(g20370) );
INV_X32 U_g20371 ( .A(g17471), .ZN(g20371) );
INV_X32 U_g20372 ( .A(g17476), .ZN(g20372) );
INV_X32 U_g20373 ( .A(g17479), .ZN(g20373) );
INV_X32 U_g20374 ( .A(g17482), .ZN(g20374) );
INV_X32 U_I26796 ( .A(g17224), .ZN(I26796) );
INV_X32 U_g20377 ( .A(I26796), .ZN(g20377) );
INV_X32 U_g20378 ( .A(g17487), .ZN(g20378) );
INV_X32 U_g20379 ( .A(g17490), .ZN(g20379) );
INV_X32 U_g20380 ( .A(g17493), .ZN(g20380) );
INV_X32 U_g20381 ( .A(g17496), .ZN(g20381) );
INV_X32 U_g20382 ( .A(g17500), .ZN(g20382) );
INV_X32 U_g20383 ( .A(g17503), .ZN(g20383) );
INV_X32 U_g20384 ( .A(g17511), .ZN(g20384) );
INV_X32 U_g20385 ( .A(g17514), .ZN(g20385) );
INV_X32 U_g20386 ( .A(g17517), .ZN(g20386) );
INV_X32 U_g20387 ( .A(g17520), .ZN(g20387) );
INV_X32 U_g20388 ( .A(g17523), .ZN(g20388) );
INV_X32 U_g20389 ( .A(g17531), .ZN(g20389) );
INV_X32 U_g20390 ( .A(g17534), .ZN(g20390) );
INV_X32 U_g20391 ( .A(g17537), .ZN(g20391) );
INV_X32 U_g20392 ( .A(g17545), .ZN(g20392) );
INV_X32 U_g20393 ( .A(g17548), .ZN(g20393) );
INV_X32 U_g20394 ( .A(g17551), .ZN(g20394) );
INV_X32 U_I26816 ( .A(g17225), .ZN(I26816) );
INV_X32 U_g20395 ( .A(I26816), .ZN(g20395) );
INV_X32 U_I26819 ( .A(g17226), .ZN(I26819) );
INV_X32 U_g20396 ( .A(I26819), .ZN(g20396) );
INV_X32 U_g20397 ( .A(g17557), .ZN(g20397) );
INV_X32 U_g20398 ( .A(g17560), .ZN(g20398) );
INV_X32 U_g20399 ( .A(g17563), .ZN(g20399) );
INV_X32 U_g20400 ( .A(g17567), .ZN(g20400) );
INV_X32 U_g20401 ( .A(g17570), .ZN(g20401) );
INV_X32 U_g20402 ( .A(g17573), .ZN(g20402) );
INV_X32 U_g20403 ( .A(g17579), .ZN(g20403) );
INV_X32 U_g20404 ( .A(g17582), .ZN(g20404) );
INV_X32 U_g20405 ( .A(g17585), .ZN(g20405) );
INV_X32 U_g20406 ( .A(g17588), .ZN(g20406) );
INV_X32 U_g20407 ( .A(g17591), .ZN(g20407) );
INV_X32 U_g20408 ( .A(g17594), .ZN(g20408) );
INV_X32 U_g20409 ( .A(g17601), .ZN(g20409) );
INV_X32 U_g20410 ( .A(g17604), .ZN(g20410) );
INV_X32 U_g20411 ( .A(g17607), .ZN(g20411) );
INV_X32 U_g20412 ( .A(g17610), .ZN(g20412) );
INV_X32 U_g20413 ( .A(g17613), .ZN(g20413) );
INV_X32 U_g20414 ( .A(g17621), .ZN(g20414) );
INV_X32 U_g20415 ( .A(g17624), .ZN(g20415) );
INV_X32 U_g20416 ( .A(g17627), .ZN(g20416) );
INV_X32 U_I26843 ( .A(g17228), .ZN(I26843) );
INV_X32 U_g20418 ( .A(I26843), .ZN(g20418) );
INV_X32 U_I26846 ( .A(g17229), .ZN(I26846) );
INV_X32 U_g20419 ( .A(I26846), .ZN(g20419) );
INV_X32 U_g20420 ( .A(g17637), .ZN(g20420) );
INV_X32 U_g20421 ( .A(g17649), .ZN(g20421) );
INV_X32 U_g20422 ( .A(g17655), .ZN(g20422) );
INV_X32 U_g20423 ( .A(g17658), .ZN(g20423) );
INV_X32 U_g20424 ( .A(g17661), .ZN(g20424) );
INV_X32 U_g20425 ( .A(g17664), .ZN(g20425) );
INV_X32 U_g20426 ( .A(g17667), .ZN(g20426) );
INV_X32 U_g20427 ( .A(g17670), .ZN(g20427) );
INV_X32 U_g20428 ( .A(g17676), .ZN(g20428) );
INV_X32 U_g20429 ( .A(g17679), .ZN(g20429) );
INV_X32 U_g20430 ( .A(g17682), .ZN(g20430) );
INV_X32 U_g20431 ( .A(g17685), .ZN(g20431) );
INV_X32 U_g20432 ( .A(g17688), .ZN(g20432) );
INV_X32 U_g20433 ( .A(g17691), .ZN(g20433) );
INV_X32 U_g20434 ( .A(g17698), .ZN(g20434) );
INV_X32 U_g20435 ( .A(g17701), .ZN(g20435) );
INV_X32 U_g20436 ( .A(g17704), .ZN(g20436) );
INV_X32 U_g20437 ( .A(g17707), .ZN(g20437) );
INV_X32 U_g20438 ( .A(g17710), .ZN(g20438) );
INV_X32 U_I26868 ( .A(g17234), .ZN(I26868) );
INV_X32 U_g20439 ( .A(I26868), .ZN(g20439) );
INV_X32 U_I26871 ( .A(g17235), .ZN(I26871) );
INV_X32 U_g20440 ( .A(I26871), .ZN(g20440) );
INV_X32 U_I26874 ( .A(g17236), .ZN(I26874) );
INV_X32 U_g20441 ( .A(I26874), .ZN(g20441) );
INV_X32 U_g20442 ( .A(g17738), .ZN(g20442) );
INV_X32 U_g20443 ( .A(g17749), .ZN(g20443) );
INV_X32 U_g20444 ( .A(g17755), .ZN(g20444) );
INV_X32 U_g20445 ( .A(g17758), .ZN(g20445) );
INV_X32 U_g20446 ( .A(g17761), .ZN(g20446) );
INV_X32 U_g20447 ( .A(g17764), .ZN(g20447) );
INV_X32 U_g20448 ( .A(g17767), .ZN(g20448) );
INV_X32 U_g20449 ( .A(g17770), .ZN(g20449) );
INV_X32 U_g20450 ( .A(g17776), .ZN(g20450) );
INV_X32 U_g20451 ( .A(g17779), .ZN(g20451) );
INV_X32 U_g20452 ( .A(g17782), .ZN(g20452) );
INV_X32 U_g20453 ( .A(g17785), .ZN(g20453) );
INV_X32 U_g20454 ( .A(g17788), .ZN(g20454) );
INV_X32 U_g20455 ( .A(g17791), .ZN(g20455) );
INV_X32 U_g20456 ( .A(g17799), .ZN(g20456) );
INV_X32 U_I26892 ( .A(g17246), .ZN(I26892) );
INV_X32 U_g20457 ( .A(I26892), .ZN(g20457) );
INV_X32 U_I26895 ( .A(g17247), .ZN(I26895) );
INV_X32 U_g20458 ( .A(I26895), .ZN(g20458) );
INV_X32 U_I26898 ( .A(g17248), .ZN(I26898) );
INV_X32 U_g20459 ( .A(I26898), .ZN(g20459) );
INV_X32 U_g20461 ( .A(g17839), .ZN(g20461) );
INV_X32 U_g20462 ( .A(g17850), .ZN(g20462) );
INV_X32 U_g20463 ( .A(g17856), .ZN(g20463) );
INV_X32 U_g20464 ( .A(g17859), .ZN(g20464) );
INV_X32 U_g20465 ( .A(g17862), .ZN(g20465) );
INV_X32 U_g20466 ( .A(g17865), .ZN(g20466) );
INV_X32 U_g20467 ( .A(g17868), .ZN(g20467) );
INV_X32 U_g20468 ( .A(g17871), .ZN(g20468) );
INV_X32 U_I26910 ( .A(g17269), .ZN(I26910) );
INV_X32 U_g20469 ( .A(I26910), .ZN(g20469) );
INV_X32 U_I26913 ( .A(g17270), .ZN(I26913) );
INV_X32 U_g20470 ( .A(I26913), .ZN(g20470) );
INV_X32 U_I26916 ( .A(g17271), .ZN(I26916) );
INV_X32 U_g20471 ( .A(I26916), .ZN(g20471) );
INV_X32 U_g20476 ( .A(g17951), .ZN(g20476) );
INV_X32 U_g20477 ( .A(g17962), .ZN(g20477) );
INV_X32 U_I26923 ( .A(g17302), .ZN(I26923) );
INV_X32 U_g20478 ( .A(I26923), .ZN(g20478) );
INV_X32 U_I26926 ( .A(g17303), .ZN(I26926) );
INV_X32 U_g20479 ( .A(I26926), .ZN(g20479) );
INV_X32 U_I26931 ( .A(g17340), .ZN(I26931) );
INV_X32 U_g20484 ( .A(I26931), .ZN(g20484) );
INV_X32 U_I26934 ( .A(g17341), .ZN(I26934) );
INV_X32 U_g20485 ( .A(I26934), .ZN(g20485) );
INV_X32 U_g20490 ( .A(g18166), .ZN(g20490) );
INV_X32 U_I26940 ( .A(g17383), .ZN(I26940) );
INV_X32 U_g20491 ( .A(I26940), .ZN(g20491) );
INV_X32 U_g20496 ( .A(g18258), .ZN(g20496) );
INV_X32 U_I26947 ( .A(g17429), .ZN(I26947) );
INV_X32 U_g20498 ( .A(I26947), .ZN(g20498) );
INV_X32 U_g20500 ( .A(g18278), .ZN(g20500) );
INV_X32 U_g20501 ( .A(g18334), .ZN(g20501) );
INV_X32 U_g20504 ( .A(g18355), .ZN(g20504) );
INV_X32 U_g20505 ( .A(g18371), .ZN(g20505) );
INV_X32 U_g20507 ( .A(g18351), .ZN(g20507) );
INV_X32 U_I26960 ( .A(g16884), .ZN(I26960) );
INV_X32 U_g20513 ( .A(I26960), .ZN(g20513) );
INV_X32 U_g20516 ( .A(g18432), .ZN(g20516) );
INV_X32 U_g20517 ( .A(g18450), .ZN(g20517) );
INV_X32 U_g20518 ( .A(g18466), .ZN(g20518) );
INV_X32 U_I26966 ( .A(g17051), .ZN(I26966) );
INV_X32 U_g20519 ( .A(I26966), .ZN(g20519) );
INV_X32 U_g20526 ( .A(g18446), .ZN(g20526) );
INV_X32 U_I26972 ( .A(g16913), .ZN(I26972) );
INV_X32 U_g20531 ( .A(I26972), .ZN(g20531) );
INV_X32 U_g20534 ( .A(g18505), .ZN(g20534) );
INV_X32 U_g20535 ( .A(g18523), .ZN(g20535) );
INV_X32 U_g20536 ( .A(g18539), .ZN(g20536) );
INV_X32 U_I26980 ( .A(g17086), .ZN(I26980) );
INV_X32 U_g20539 ( .A(I26980), .ZN(g20539) );
INV_X32 U_g20545 ( .A(g18519), .ZN(g20545) );
INV_X32 U_I26985 ( .A(g16943), .ZN(I26985) );
INV_X32 U_g20550 ( .A(I26985), .ZN(g20550) );
INV_X32 U_g20553 ( .A(g18569), .ZN(g20553) );
INV_X32 U_g20554 ( .A(g18587), .ZN(g20554) );
INV_X32 U_I26990 ( .A(g19145), .ZN(I26990) );
INV_X32 U_g20555 ( .A(I26990), .ZN(g20555) );
INV_X32 U_I26993 ( .A(g19159), .ZN(I26993) );
INV_X32 U_g20556 ( .A(I26993), .ZN(g20556) );
INV_X32 U_I26996 ( .A(g19169), .ZN(I26996) );
INV_X32 U_g20557 ( .A(I26996), .ZN(g20557) );
INV_X32 U_I26999 ( .A(g19543), .ZN(I26999) );
INV_X32 U_g20558 ( .A(I26999), .ZN(g20558) );
INV_X32 U_I27002 ( .A(g19147), .ZN(I27002) );
INV_X32 U_g20559 ( .A(I27002), .ZN(g20559) );
INV_X32 U_I27005 ( .A(g19164), .ZN(I27005) );
INV_X32 U_g20560 ( .A(I27005), .ZN(g20560) );
INV_X32 U_I27008 ( .A(g19175), .ZN(I27008) );
INV_X32 U_g20561 ( .A(I27008), .ZN(g20561) );
INV_X32 U_I27011 ( .A(g19546), .ZN(I27011) );
INV_X32 U_g20562 ( .A(I27011), .ZN(g20562) );
INV_X32 U_I27014 ( .A(g19151), .ZN(I27014) );
INV_X32 U_g20563 ( .A(I27014), .ZN(g20563) );
INV_X32 U_I27017 ( .A(g19170), .ZN(I27017) );
INV_X32 U_g20564 ( .A(I27017), .ZN(g20564) );
INV_X32 U_I27020 ( .A(g19182), .ZN(I27020) );
INV_X32 U_g20565 ( .A(I27020), .ZN(g20565) );
INV_X32 U_I27023 ( .A(g19550), .ZN(I27023) );
INV_X32 U_g20566 ( .A(I27023), .ZN(g20566) );
INV_X32 U_I27026 ( .A(g19156), .ZN(I27026) );
INV_X32 U_g20567 ( .A(I27026), .ZN(g20567) );
INV_X32 U_I27029 ( .A(g19176), .ZN(I27029) );
INV_X32 U_g20568 ( .A(I27029), .ZN(g20568) );
INV_X32 U_I27032 ( .A(g19189), .ZN(I27032) );
INV_X32 U_g20569 ( .A(I27032), .ZN(g20569) );
INV_X32 U_I27035 ( .A(g19556), .ZN(I27035) );
INV_X32 U_g20570 ( .A(I27035), .ZN(g20570) );
INV_X32 U_I27038 ( .A(g20082), .ZN(I27038) );
INV_X32 U_g20571 ( .A(I27038), .ZN(g20571) );
INV_X32 U_I27041 ( .A(g19237), .ZN(I27041) );
INV_X32 U_g20572 ( .A(I27041), .ZN(g20572) );
INV_X32 U_I27044 ( .A(g19247), .ZN(I27044) );
INV_X32 U_g20573 ( .A(I27044), .ZN(g20573) );
INV_X32 U_I27047 ( .A(g19258), .ZN(I27047) );
INV_X32 U_g20574 ( .A(I27047), .ZN(g20574) );
INV_X32 U_I27050 ( .A(g19183), .ZN(I27050) );
INV_X32 U_g20575 ( .A(I27050), .ZN(g20575) );
INV_X32 U_I27053 ( .A(g19190), .ZN(I27053) );
INV_X32 U_g20576 ( .A(I27053), .ZN(g20576) );
INV_X32 U_I27056 ( .A(g19196), .ZN(I27056) );
INV_X32 U_g20577 ( .A(I27056), .ZN(g20577) );
INV_X32 U_I27059 ( .A(g19207), .ZN(I27059) );
INV_X32 U_g20578 ( .A(I27059), .ZN(g20578) );
INV_X32 U_I27062 ( .A(g19217), .ZN(I27062) );
INV_X32 U_g20579 ( .A(I27062), .ZN(g20579) );
INV_X32 U_I27065 ( .A(g19270), .ZN(I27065) );
INV_X32 U_g20580 ( .A(I27065), .ZN(g20580) );
INV_X32 U_I27068 ( .A(g19197), .ZN(I27068) );
INV_X32 U_g20581 ( .A(I27068), .ZN(g20581) );
INV_X32 U_I27071 ( .A(g19218), .ZN(I27071) );
INV_X32 U_g20582 ( .A(I27071), .ZN(g20582) );
INV_X32 U_I27074 ( .A(g19238), .ZN(I27074) );
INV_X32 U_g20583 ( .A(I27074), .ZN(g20583) );
INV_X32 U_I27077 ( .A(g19259), .ZN(I27077) );
INV_X32 U_g20584 ( .A(I27077), .ZN(g20584) );
INV_X32 U_I27080 ( .A(g19198), .ZN(I27080) );
INV_X32 U_g20585 ( .A(I27080), .ZN(g20585) );
INV_X32 U_I27083 ( .A(g19208), .ZN(I27083) );
INV_X32 U_g20586 ( .A(I27083), .ZN(g20586) );
INV_X32 U_I27086 ( .A(g19229), .ZN(I27086) );
INV_X32 U_g20587 ( .A(I27086), .ZN(g20587) );
INV_X32 U_I27089 ( .A(g20105), .ZN(I27089) );
INV_X32 U_g20588 ( .A(I27089), .ZN(g20588) );
INV_X32 U_I27092 ( .A(g19174), .ZN(I27092) );
INV_X32 U_g20589 ( .A(I27092), .ZN(g20589) );
INV_X32 U_I27095 ( .A(g19185), .ZN(I27095) );
INV_X32 U_g20590 ( .A(I27095), .ZN(g20590) );
INV_X32 U_I27098 ( .A(g19199), .ZN(I27098) );
INV_X32 U_g20591 ( .A(I27098), .ZN(g20591) );
INV_X32 U_I27101 ( .A(g19220), .ZN(I27101) );
INV_X32 U_g20592 ( .A(I27101), .ZN(g20592) );
INV_X32 U_I27104 ( .A(g19239), .ZN(I27104) );
INV_X32 U_g20593 ( .A(I27104), .ZN(g20593) );
INV_X32 U_I27107 ( .A(g19249), .ZN(I27107) );
INV_X32 U_g20594 ( .A(I27107), .ZN(g20594) );
INV_X32 U_I27110 ( .A(g19622), .ZN(I27110) );
INV_X32 U_g20595 ( .A(I27110), .ZN(g20595) );
INV_X32 U_I27113 ( .A(g19689), .ZN(I27113) );
INV_X32 U_g20596 ( .A(I27113), .ZN(g20596) );
INV_X32 U_I27116 ( .A(g19762), .ZN(I27116) );
INV_X32 U_g20597 ( .A(I27116), .ZN(g20597) );
INV_X32 U_I27119 ( .A(g19563), .ZN(I27119) );
INV_X32 U_g20598 ( .A(I27119), .ZN(g20598) );
INV_X32 U_I27122 ( .A(g19595), .ZN(I27122) );
INV_X32 U_g20599 ( .A(I27122), .ZN(g20599) );
INV_X32 U_I27125 ( .A(g19652), .ZN(I27125) );
INV_X32 U_g20600 ( .A(I27125), .ZN(g20600) );
INV_X32 U_I27128 ( .A(g19725), .ZN(I27128) );
INV_X32 U_g20601 ( .A(I27128), .ZN(g20601) );
INV_X32 U_I27131 ( .A(g19798), .ZN(I27131) );
INV_X32 U_g20602 ( .A(I27131), .ZN(g20602) );
INV_X32 U_I27134 ( .A(g19573), .ZN(I27134) );
INV_X32 U_g20603 ( .A(I27134), .ZN(g20603) );
INV_X32 U_I27137 ( .A(g19596), .ZN(I27137) );
INV_X32 U_g20604 ( .A(I27137), .ZN(g20604) );
INV_X32 U_I27140 ( .A(g19690), .ZN(I27140) );
INV_X32 U_g20605 ( .A(I27140), .ZN(g20605) );
INV_X32 U_I27143 ( .A(g19763), .ZN(I27143) );
INV_X32 U_g20606 ( .A(I27143), .ZN(g20606) );
INV_X32 U_I27146 ( .A(g19838), .ZN(I27146) );
INV_X32 U_g20607 ( .A(I27146), .ZN(g20607) );
INV_X32 U_I27149 ( .A(g19893), .ZN(I27149) );
INV_X32 U_g20608 ( .A(I27149), .ZN(g20608) );
INV_X32 U_I27152 ( .A(g20360), .ZN(I27152) );
INV_X32 U_g20609 ( .A(I27152), .ZN(g20609) );
INV_X32 U_I27155 ( .A(g20395), .ZN(I27155) );
INV_X32 U_g20610 ( .A(I27155), .ZN(g20610) );
INV_X32 U_I27158 ( .A(g20439), .ZN(I27158) );
INV_X32 U_g20611 ( .A(I27158), .ZN(g20611) );
INV_X32 U_I27161 ( .A(g20377), .ZN(I27161) );
INV_X32 U_g20612 ( .A(I27161), .ZN(g20612) );
INV_X32 U_I27164 ( .A(g20418), .ZN(I27164) );
INV_X32 U_g20613 ( .A(I27164), .ZN(g20613) );
INV_X32 U_I27167 ( .A(g20457), .ZN(I27167) );
INV_X32 U_g20614 ( .A(I27167), .ZN(g20614) );
INV_X32 U_I27170 ( .A(g20396), .ZN(I27170) );
INV_X32 U_g20615 ( .A(I27170), .ZN(g20615) );
INV_X32 U_I27173 ( .A(g20440), .ZN(I27173) );
INV_X32 U_g20616 ( .A(I27173), .ZN(g20616) );
INV_X32 U_I27176 ( .A(g20469), .ZN(I27176) );
INV_X32 U_g20617 ( .A(I27176), .ZN(g20617) );
INV_X32 U_I27179 ( .A(g20419), .ZN(I27179) );
INV_X32 U_g20618 ( .A(I27179), .ZN(g20618) );
INV_X32 U_I27182 ( .A(g20458), .ZN(I27182) );
INV_X32 U_g20619 ( .A(I27182), .ZN(g20619) );
INV_X32 U_I27185 ( .A(g20478), .ZN(I27185) );
INV_X32 U_g20620 ( .A(I27185), .ZN(g20620) );
INV_X32 U_I27188 ( .A(g20441), .ZN(I27188) );
INV_X32 U_g20621 ( .A(I27188), .ZN(g20621) );
INV_X32 U_I27191 ( .A(g20470), .ZN(I27191) );
INV_X32 U_g20622 ( .A(I27191), .ZN(g20622) );
INV_X32 U_I27194 ( .A(g20484), .ZN(I27194) );
INV_X32 U_g20623 ( .A(I27194), .ZN(g20623) );
INV_X32 U_I27197 ( .A(g20459), .ZN(I27197) );
INV_X32 U_g20624 ( .A(I27197), .ZN(g20624) );
INV_X32 U_I27200 ( .A(g20479), .ZN(I27200) );
INV_X32 U_g20625 ( .A(I27200), .ZN(g20625) );
INV_X32 U_I27203 ( .A(g20491), .ZN(I27203) );
INV_X32 U_g20626 ( .A(I27203), .ZN(g20626) );
INV_X32 U_I27206 ( .A(g20471), .ZN(I27206) );
INV_X32 U_g20627 ( .A(I27206), .ZN(g20627) );
INV_X32 U_I27209 ( .A(g20485), .ZN(I27209) );
INV_X32 U_g20628 ( .A(I27209), .ZN(g20628) );
INV_X32 U_I27212 ( .A(g20498), .ZN(I27212) );
INV_X32 U_g20629 ( .A(I27212), .ZN(g20629) );
INV_X32 U_I27215 ( .A(g19158), .ZN(I27215) );
INV_X32 U_g20630 ( .A(I27215), .ZN(g20630) );
INV_X32 U_I27218 ( .A(g19168), .ZN(I27218) );
INV_X32 U_g20631 ( .A(I27218), .ZN(g20631) );
INV_X32 U_I27221 ( .A(g19180), .ZN(I27221) );
INV_X32 U_g20632 ( .A(I27221), .ZN(g20632) );
INV_X32 U_I27225 ( .A(g19358), .ZN(I27225) );
INV_X32 U_g20634 ( .A(I27225), .ZN(g20634) );
INV_X32 U_I27228 ( .A(g19390), .ZN(I27228) );
INV_X32 U_g20637 ( .A(I27228), .ZN(g20637) );
INV_X32 U_I27232 ( .A(g19401), .ZN(I27232) );
INV_X32 U_g20641 ( .A(I27232), .ZN(g20641) );
INV_X32 U_I27235 ( .A(g19420), .ZN(I27235) );
INV_X32 U_g20644 ( .A(I27235), .ZN(g20644) );
INV_X32 U_I27240 ( .A(g19335), .ZN(I27240) );
INV_X32 U_g20649 ( .A(I27240), .ZN(g20649) );
INV_X32 U_I27243 ( .A(g19335), .ZN(I27243) );
INV_X32 U_g20652 ( .A(I27243), .ZN(g20652) );
INV_X32 U_I27246 ( .A(g19335), .ZN(I27246) );
INV_X32 U_g20655 ( .A(I27246), .ZN(g20655) );
INV_X32 U_I27250 ( .A(g19390), .ZN(I27250) );
INV_X32 U_g20659 ( .A(I27250), .ZN(g20659) );
INV_X32 U_I27253 ( .A(g19420), .ZN(I27253) );
INV_X32 U_g20662 ( .A(I27253), .ZN(g20662) );
INV_X32 U_I27257 ( .A(g19431), .ZN(I27257) );
INV_X32 U_g20666 ( .A(I27257), .ZN(g20666) );
INV_X32 U_I27260 ( .A(g19457), .ZN(I27260) );
INV_X32 U_g20669 ( .A(I27260), .ZN(g20669) );
INV_X32 U_I27264 ( .A(g19358), .ZN(I27264) );
INV_X32 U_g20673 ( .A(I27264), .ZN(g20673) );
INV_X32 U_I27267 ( .A(g19358), .ZN(I27267) );
INV_X32 U_g20676 ( .A(I27267), .ZN(g20676) );
INV_X32 U_I27270 ( .A(g19335), .ZN(I27270) );
INV_X32 U_g20679 ( .A(I27270), .ZN(g20679) );
INV_X32 U_I27275 ( .A(g19369), .ZN(I27275) );
INV_X32 U_g20684 ( .A(I27275), .ZN(g20684) );
INV_X32 U_I27278 ( .A(g19369), .ZN(I27278) );
INV_X32 U_g20687 ( .A(I27278), .ZN(g20687) );
INV_X32 U_I27281 ( .A(g19369), .ZN(I27281) );
INV_X32 U_g20690 ( .A(I27281), .ZN(g20690) );
INV_X32 U_I27285 ( .A(g19420), .ZN(I27285) );
INV_X32 U_g20694 ( .A(I27285), .ZN(g20694) );
INV_X32 U_I27288 ( .A(g19457), .ZN(I27288) );
INV_X32 U_g20697 ( .A(I27288), .ZN(g20697) );
INV_X32 U_I27293 ( .A(g19335), .ZN(I27293) );
INV_X32 U_g20704 ( .A(I27293), .ZN(g20704) );
INV_X32 U_I27297 ( .A(g19390), .ZN(I27297) );
INV_X32 U_g20708 ( .A(I27297), .ZN(g20708) );
INV_X32 U_I27300 ( .A(g19390), .ZN(I27300) );
INV_X32 U_g20711 ( .A(I27300), .ZN(g20711) );
INV_X32 U_I27303 ( .A(g19369), .ZN(I27303) );
INV_X32 U_g20714 ( .A(I27303), .ZN(g20714) );
INV_X32 U_I27308 ( .A(g19401), .ZN(I27308) );
INV_X32 U_g20719 ( .A(I27308), .ZN(g20719) );
INV_X32 U_I27311 ( .A(g19401), .ZN(I27311) );
INV_X32 U_g20722 ( .A(I27311), .ZN(g20722) );
INV_X32 U_I27314 ( .A(g19401), .ZN(I27314) );
INV_X32 U_g20725 ( .A(I27314), .ZN(g20725) );
INV_X32 U_I27318 ( .A(g19457), .ZN(I27318) );
INV_X32 U_g20729 ( .A(I27318), .ZN(g20729) );
INV_X32 U_I27321 ( .A(g19335), .ZN(I27321) );
INV_X32 U_g20732 ( .A(I27321), .ZN(g20732) );
INV_X32 U_I27324 ( .A(g19358), .ZN(I27324) );
INV_X32 U_g20735 ( .A(I27324), .ZN(g20735) );
INV_X32 U_I27328 ( .A(g19369), .ZN(I27328) );
INV_X32 U_g20739 ( .A(I27328), .ZN(g20739) );
INV_X32 U_I27332 ( .A(g19420), .ZN(I27332) );
INV_X32 U_g20743 ( .A(I27332), .ZN(g20743) );
INV_X32 U_I27335 ( .A(g19420), .ZN(I27335) );
INV_X32 U_g20746 ( .A(I27335), .ZN(g20746) );
INV_X32 U_I27338 ( .A(g19401), .ZN(I27338) );
INV_X32 U_g20749 ( .A(I27338), .ZN(g20749) );
INV_X32 U_I27343 ( .A(g19431), .ZN(I27343) );
INV_X32 U_g20754 ( .A(I27343), .ZN(g20754) );
INV_X32 U_I27346 ( .A(g19431), .ZN(I27346) );
INV_X32 U_g20757 ( .A(I27346), .ZN(g20757) );
INV_X32 U_I27349 ( .A(g19431), .ZN(I27349) );
INV_X32 U_g20760 ( .A(I27349), .ZN(g20760) );
INV_X32 U_I27352 ( .A(g19358), .ZN(I27352) );
INV_X32 U_g20763 ( .A(I27352), .ZN(g20763) );
INV_X32 U_I27355 ( .A(g19335), .ZN(I27355) );
INV_X32 U_g20766 ( .A(I27355), .ZN(g20766) );
INV_X32 U_I27358 ( .A(g19369), .ZN(I27358) );
INV_X32 U_g20769 ( .A(I27358), .ZN(g20769) );
INV_X32 U_I27361 ( .A(g19390), .ZN(I27361) );
INV_X32 U_g20772 ( .A(I27361), .ZN(g20772) );
INV_X32 U_I27365 ( .A(g19401), .ZN(I27365) );
INV_X32 U_g20776 ( .A(I27365), .ZN(g20776) );
INV_X32 U_I27369 ( .A(g19457), .ZN(I27369) );
INV_X32 U_g20780 ( .A(I27369), .ZN(g20780) );
INV_X32 U_I27372 ( .A(g19457), .ZN(I27372) );
INV_X32 U_g20783 ( .A(I27372), .ZN(g20783) );
INV_X32 U_I27375 ( .A(g19431), .ZN(I27375) );
INV_X32 U_g20786 ( .A(I27375), .ZN(g20786) );
INV_X32 U_I27379 ( .A(g19358), .ZN(I27379) );
INV_X32 U_g20790 ( .A(I27379), .ZN(g20790) );
INV_X32 U_I27382 ( .A(g19390), .ZN(I27382) );
INV_X32 U_g20793 ( .A(I27382), .ZN(g20793) );
INV_X32 U_I27385 ( .A(g19369), .ZN(I27385) );
INV_X32 U_g20796 ( .A(I27385), .ZN(g20796) );
INV_X32 U_I27388 ( .A(g19401), .ZN(I27388) );
INV_X32 U_g20799 ( .A(I27388), .ZN(g20799) );
INV_X32 U_I27391 ( .A(g19420), .ZN(I27391) );
INV_X32 U_g20802 ( .A(I27391), .ZN(g20802) );
INV_X32 U_I27395 ( .A(g19431), .ZN(I27395) );
INV_X32 U_g20806 ( .A(I27395), .ZN(g20806) );
INV_X32 U_I27399 ( .A(g19390), .ZN(I27399) );
INV_X32 U_g20810 ( .A(I27399), .ZN(g20810) );
INV_X32 U_I27402 ( .A(g19420), .ZN(I27402) );
INV_X32 U_g20813 ( .A(I27402), .ZN(g20813) );
INV_X32 U_I27405 ( .A(g19401), .ZN(I27405) );
INV_X32 U_g20816 ( .A(I27405), .ZN(g20816) );
INV_X32 U_I27408 ( .A(g19431), .ZN(I27408) );
INV_X32 U_g20819 ( .A(I27408), .ZN(g20819) );
INV_X32 U_I27411 ( .A(g19457), .ZN(I27411) );
INV_X32 U_g20822 ( .A(I27411), .ZN(g20822) );
INV_X32 U_I27416 ( .A(g19420), .ZN(I27416) );
INV_X32 U_g20827 ( .A(I27416), .ZN(g20827) );
INV_X32 U_I27419 ( .A(g19457), .ZN(I27419) );
INV_X32 U_g20830 ( .A(I27419), .ZN(g20830) );
INV_X32 U_I27422 ( .A(g19431), .ZN(I27422) );
INV_X32 U_g20833 ( .A(I27422), .ZN(g20833) );
INV_X32 U_I27426 ( .A(g19457), .ZN(I27426) );
INV_X32 U_g20837 ( .A(I27426), .ZN(g20837) );
INV_X32 U_g20842 ( .A(g19441), .ZN(g20842) );
INV_X32 U_g20850 ( .A(g19468), .ZN(g20850) );
INV_X32 U_g20858 ( .A(g19491), .ZN(g20858) );
INV_X32 U_g20866 ( .A(g19512), .ZN(g20866) );
INV_X32 U_g20885 ( .A(g19865), .ZN(g20885) );
INV_X32 U_g20904 ( .A(g19896), .ZN(g20904) );
INV_X32 U_g20928 ( .A(g19921), .ZN(g20928) );
INV_X32 U_I27488 ( .A(g20310), .ZN(I27488) );
INV_X32 U_g20942 ( .A(I27488), .ZN(g20942) );
INV_X32 U_I27491 ( .A(g20314), .ZN(I27491) );
INV_X32 U_g20943 ( .A(I27491), .ZN(g20943) );
INV_X32 U_g20956 ( .A(g19936), .ZN(g20956) );
INV_X32 U_I27516 ( .A(g20333), .ZN(I27516) );
INV_X32 U_g20971 ( .A(I27516), .ZN(g20971) );
INV_X32 U_I27531 ( .A(g20343), .ZN(I27531) );
INV_X32 U_g20984 ( .A(I27531), .ZN(g20984) );
INV_X32 U_I27534 ( .A(g20083), .ZN(I27534) );
INV_X32 U_g20985 ( .A(I27534), .ZN(g20985) );
INV_X32 U_I27537 ( .A(g19957), .ZN(I27537) );
INV_X32 U_g20986 ( .A(I27537), .ZN(g20986) );
INV_X32 U_I27549 ( .A(g20353), .ZN(I27549) );
INV_X32 U_g20998 ( .A(I27549), .ZN(g20998) );
INV_X32 U_I27565 ( .A(g19987), .ZN(I27565) );
INV_X32 U_g21012 ( .A(I27565), .ZN(g21012) );
INV_X32 U_I27577 ( .A(g20375), .ZN(I27577) );
INV_X32 U_g21024 ( .A(I27577), .ZN(g21024) );
INV_X32 U_I27585 ( .A(g20376), .ZN(I27585) );
INV_X32 U_g21030 ( .A(I27585), .ZN(g21030) );
INV_X32 U_I27593 ( .A(g20025), .ZN(I27593) );
INV_X32 U_g21036 ( .A(I27593), .ZN(g21036) );
INV_X32 U_g21050 ( .A(g20513), .ZN(g21050) );
INV_X32 U_I27614 ( .A(g20067), .ZN(I27614) );
INV_X32 U_g21057 ( .A(I27614), .ZN(g21057) );
INV_X32 U_I27621 ( .A(g20417), .ZN(I27621) );
INV_X32 U_g21064 ( .A(I27621), .ZN(g21064) );
INV_X32 U_g21066 ( .A(g20519), .ZN(g21066) );
INV_X32 U_g21069 ( .A(g20531), .ZN(g21069) );
INV_X32 U_g21076 ( .A(g20539), .ZN(g21076) );
INV_X32 U_g21079 ( .A(g20550), .ZN(g21079) );
INV_X32 U_I27646 ( .A(g20507), .ZN(I27646) );
INV_X32 U_g21087 ( .A(I27646), .ZN(g21087) );
INV_X32 U_g21090 ( .A(g19064), .ZN(g21090) );
INV_X32 U_g21093 ( .A(g19075), .ZN(g21093) );
INV_X32 U_I27658 ( .A(g20526), .ZN(I27658) );
INV_X32 U_g21099 ( .A(I27658), .ZN(g21099) );
INV_X32 U_g21102 ( .A(g19081), .ZN(g21102) );
INV_X32 U_I27667 ( .A(g20507), .ZN(I27667) );
INV_X32 U_g21108 ( .A(I27667), .ZN(g21108) );
INV_X32 U_I27672 ( .A(g20545), .ZN(I27672) );
INV_X32 U_g21113 ( .A(I27672), .ZN(g21113) );
INV_X32 U_I27684 ( .A(g20526), .ZN(I27684) );
INV_X32 U_g21125 ( .A(I27684), .ZN(g21125) );
INV_X32 U_I27689 ( .A(g19070), .ZN(I27689) );
INV_X32 U_g21130 ( .A(I27689), .ZN(g21130) );
INV_X32 U_I27705 ( .A(g20545), .ZN(I27705) );
INV_X32 U_g21144 ( .A(I27705), .ZN(g21144) );
INV_X32 U_I27727 ( .A(g19070), .ZN(I27727) );
INV_X32 U_g21164 ( .A(I27727), .ZN(g21164) );
INV_X32 U_I27749 ( .A(g19954), .ZN(I27749) );
INV_X32 U_g21184 ( .A(I27749), .ZN(g21184) );
INV_X32 U_g21187 ( .A(g19113), .ZN(g21187) );
INV_X32 U_I27766 ( .A(g19984), .ZN(I27766) );
INV_X32 U_g21199 ( .A(I27766), .ZN(g21199) );
INV_X32 U_g21202 ( .A(g19118), .ZN(g21202) );
INV_X32 U_I27779 ( .A(g20022), .ZN(I27779) );
INV_X32 U_g21214 ( .A(I27779), .ZN(g21214) );
INV_X32 U_g21217 ( .A(g19125), .ZN(g21217) );
INV_X32 U_I27785 ( .A(g20064), .ZN(I27785) );
INV_X32 U_g21222 ( .A(I27785), .ZN(g21222) );
INV_X32 U_g21225 ( .A(g19132), .ZN(g21225) );
INV_X32 U_g21241 ( .A(g19945), .ZN(g21241) );
INV_X32 U_g21249 ( .A(g19972), .ZN(g21249) );
INV_X32 U_g21258 ( .A(g20002), .ZN(g21258) );
INV_X32 U_g21266 ( .A(g20040), .ZN(g21266) );
INV_X32 U_I27822 ( .A(g19865), .ZN(I27822) );
INV_X32 U_g21271 ( .A(I27822), .ZN(g21271) );
INV_X32 U_I27827 ( .A(g19896), .ZN(I27827) );
INV_X32 U_g21278 ( .A(I27827), .ZN(g21278) );
INV_X32 U_I27832 ( .A(g19921), .ZN(I27832) );
INV_X32 U_g21285 ( .A(I27832), .ZN(g21285) );
INV_X32 U_I27838 ( .A(g19936), .ZN(I27838) );
INV_X32 U_g21293 ( .A(I27838), .ZN(g21293) );
INV_X32 U_I27868 ( .A(g19144), .ZN(I27868) );
INV_X32 U_g21327 ( .A(I27868), .ZN(g21327) );
INV_X32 U_I27897 ( .A(g19149), .ZN(I27897) );
INV_X32 U_g21358 ( .A(I27897), .ZN(g21358) );
INV_X32 U_I27900 ( .A(g19096), .ZN(I27900) );
INV_X32 U_g21359 ( .A(I27900), .ZN(g21359) );
INV_X32 U_I27917 ( .A(g19153), .ZN(I27917) );
INV_X32 U_g21376 ( .A(I27917), .ZN(g21376) );
INV_X32 U_I27920 ( .A(g19154), .ZN(I27920) );
INV_X32 U_g21377 ( .A(I27920), .ZN(g21377) );
INV_X32 U_I27927 ( .A(g19957), .ZN(I27927) );
INV_X32 U_g21382 ( .A(I27927), .ZN(g21382) );
INV_X32 U_I27942 ( .A(g19157), .ZN(I27942) );
INV_X32 U_g21399 ( .A(I27942), .ZN(g21399) );
INV_X32 U_g21400 ( .A(g19918), .ZN(g21400) );
INV_X32 U_I27949 ( .A(g19957), .ZN(I27949) );
INV_X32 U_g21404 ( .A(I27949), .ZN(g21404) );
INV_X32 U_I27958 ( .A(g19987), .ZN(I27958) );
INV_X32 U_g21415 ( .A(I27958), .ZN(g21415) );
INV_X32 U_I27969 ( .A(g19162), .ZN(I27969) );
INV_X32 U_g21426 ( .A(I27969), .ZN(g21426) );
INV_X32 U_I27972 ( .A(g19163), .ZN(I27972) );
INV_X32 U_g21427 ( .A(I27972), .ZN(g21427) );
INV_X32 U_I27976 ( .A(g19957), .ZN(I27976) );
INV_X32 U_g21429 ( .A(I27976), .ZN(g21429) );
INV_X32 U_I27984 ( .A(g19987), .ZN(I27984) );
INV_X32 U_g21441 ( .A(I27984), .ZN(g21441) );
INV_X32 U_I27992 ( .A(g20025), .ZN(I27992) );
INV_X32 U_g21449 ( .A(I27992), .ZN(g21449) );
INV_X32 U_I28000 ( .A(g19167), .ZN(I28000) );
INV_X32 U_g21457 ( .A(I28000), .ZN(g21457) );
INV_X32 U_I28003 ( .A(g19957), .ZN(I28003) );
INV_X32 U_g21458 ( .A(I28003), .ZN(g21458) );
INV_X32 U_g21461 ( .A(g19957), .ZN(g21461) );
INV_X32 U_I28009 ( .A(g20473), .ZN(I28009) );
INV_X32 U_g21473 ( .A(I28009), .ZN(g21473) );
INV_X32 U_I28013 ( .A(g19987), .ZN(I28013) );
INV_X32 U_g21477 ( .A(I28013), .ZN(g21477) );
INV_X32 U_I28019 ( .A(g20025), .ZN(I28019) );
INV_X32 U_g21483 ( .A(I28019), .ZN(g21483) );
INV_X32 U_I28027 ( .A(g20067), .ZN(I28027) );
INV_X32 U_g21491 ( .A(I28027), .ZN(g21491) );
INV_X32 U_I28031 ( .A(g19172), .ZN(I28031) );
INV_X32 U_g21495 ( .A(I28031), .ZN(g21495) );
INV_X32 U_I28034 ( .A(g19173), .ZN(I28034) );
INV_X32 U_g21496 ( .A(I28034), .ZN(g21496) );
INV_X32 U_I28038 ( .A(g19957), .ZN(I28038) );
INV_X32 U_g21498 ( .A(I28038), .ZN(g21498) );
INV_X32 U_I28043 ( .A(g19987), .ZN(I28043) );
INV_X32 U_g21505 ( .A(I28043), .ZN(g21505) );
INV_X32 U_g21508 ( .A(g19987), .ZN(g21508) );
INV_X32 U_I28047 ( .A(g20481), .ZN(I28047) );
INV_X32 U_g21514 ( .A(I28047), .ZN(g21514) );
INV_X32 U_I28051 ( .A(g20025), .ZN(I28051) );
INV_X32 U_g21518 ( .A(I28051), .ZN(g21518) );
INV_X32 U_I28057 ( .A(g20067), .ZN(I28057) );
INV_X32 U_g21524 ( .A(I28057), .ZN(g21524) );
INV_X32 U_I28061 ( .A(g19178), .ZN(I28061) );
INV_X32 U_g21528 ( .A(I28061), .ZN(g21528) );
INV_X32 U_g21529 ( .A(g19272), .ZN(g21529) );
INV_X32 U_I28065 ( .A(g19957), .ZN(I28065) );
INV_X32 U_g21530 ( .A(I28065), .ZN(g21530) );
INV_X32 U_I28072 ( .A(g19987), .ZN(I28072) );
INV_X32 U_g21537 ( .A(I28072), .ZN(g21537) );
INV_X32 U_I28076 ( .A(g20025), .ZN(I28076) );
INV_X32 U_g21541 ( .A(I28076), .ZN(g21541) );
INV_X32 U_g21544 ( .A(g20025), .ZN(g21544) );
INV_X32 U_I28080 ( .A(g20487), .ZN(I28080) );
INV_X32 U_g21550 ( .A(I28080), .ZN(g21550) );
INV_X32 U_I28084 ( .A(g20067), .ZN(I28084) );
INV_X32 U_g21554 ( .A(I28084), .ZN(g21554) );
INV_X32 U_I28087 ( .A(g19184), .ZN(I28087) );
INV_X32 U_g21557 ( .A(I28087), .ZN(g21557) );
INV_X32 U_I28090 ( .A(g20008), .ZN(I28090) );
INV_X32 U_g21558 ( .A(I28090), .ZN(g21558) );
INV_X32 U_I28093 ( .A(g19957), .ZN(I28093) );
INV_X32 U_g21561 ( .A(I28093), .ZN(g21561) );
INV_X32 U_g21565 ( .A(g19291), .ZN(g21565) );
INV_X32 U_I28100 ( .A(g19987), .ZN(I28100) );
INV_X32 U_g21566 ( .A(I28100), .ZN(g21566) );
INV_X32 U_I28107 ( .A(g20025), .ZN(I28107) );
INV_X32 U_g21573 ( .A(I28107), .ZN(g21573) );
INV_X32 U_I28111 ( .A(g20067), .ZN(I28111) );
INV_X32 U_g21577 ( .A(I28111), .ZN(g21577) );
INV_X32 U_g21580 ( .A(g20067), .ZN(g21580) );
INV_X32 U_I28115 ( .A(g20493), .ZN(I28115) );
INV_X32 U_g21586 ( .A(I28115), .ZN(g21586) );
INV_X32 U_I28119 ( .A(g19957), .ZN(I28119) );
INV_X32 U_g21590 ( .A(I28119), .ZN(g21590) );
INV_X32 U_I28123 ( .A(g19987), .ZN(I28123) );
INV_X32 U_g21594 ( .A(I28123), .ZN(g21594) );
INV_X32 U_g21598 ( .A(g19309), .ZN(g21598) );
INV_X32 U_I28130 ( .A(g20025), .ZN(I28130) );
INV_X32 U_g21599 ( .A(I28130), .ZN(g21599) );
INV_X32 U_I28137 ( .A(g20067), .ZN(I28137) );
INV_X32 U_g21606 ( .A(I28137), .ZN(g21606) );
INV_X32 U_I28143 ( .A(g19957), .ZN(I28143) );
INV_X32 U_g21612 ( .A(I28143), .ZN(g21612) );
INV_X32 U_I28148 ( .A(g19987), .ZN(I28148) );
INV_X32 U_g21619 ( .A(I28148), .ZN(g21619) );
INV_X32 U_I28152 ( .A(g20025), .ZN(I28152) );
INV_X32 U_g21623 ( .A(I28152), .ZN(g21623) );
INV_X32 U_g21627 ( .A(g19330), .ZN(g21627) );
INV_X32 U_I28159 ( .A(g20067), .ZN(I28159) );
INV_X32 U_g21628 ( .A(I28159), .ZN(g21628) );
INV_X32 U_I28169 ( .A(g19987), .ZN(I28169) );
INV_X32 U_g21640 ( .A(I28169), .ZN(g21640) );
INV_X32 U_I28174 ( .A(g20025), .ZN(I28174) );
INV_X32 U_g21647 ( .A(I28174), .ZN(g21647) );
INV_X32 U_I28178 ( .A(g20067), .ZN(I28178) );
INV_X32 U_g21651 ( .A(I28178), .ZN(g21651) );
INV_X32 U_I28184 ( .A(g19103), .ZN(I28184) );
INV_X32 U_g21655 ( .A(I28184), .ZN(g21655) );
INV_X32 U_g21661 ( .A(g19091), .ZN(g21661) );
INV_X32 U_I28201 ( .A(g20025), .ZN(I28201) );
INV_X32 U_g21671 ( .A(I28201), .ZN(g21671) );
INV_X32 U_I28206 ( .A(g20067), .ZN(I28206) );
INV_X32 U_g21678 ( .A(I28206), .ZN(g21678) );
INV_X32 U_I28210 ( .A(g20537), .ZN(I28210) );
INV_X32 U_g21682 ( .A(I28210), .ZN(g21682) );
INV_X32 U_g21690 ( .A(g19098), .ZN(g21690) );
INV_X32 U_I28229 ( .A(g20067), .ZN(I28229) );
INV_X32 U_g21700 ( .A(I28229), .ZN(g21700) );
INV_X32 U_I28235 ( .A(g20153), .ZN(I28235) );
INV_X32 U_g21708 ( .A(I28235), .ZN(g21708) );
INV_X32 U_g21716 ( .A(g19894), .ZN(g21716) );
INV_X32 U_g21726 ( .A(g19105), .ZN(g21726) );
INV_X32 U_g21742 ( .A(g19919), .ZN(g21742) );
INV_X32 U_g21752 ( .A(g19110), .ZN(g21752) );
INV_X32 U_g21766 ( .A(g19934), .ZN(g21766) );
INV_X32 U_g21782 ( .A(g19951), .ZN(g21782) );
INV_X32 U_I28314 ( .A(g19152), .ZN(I28314) );
INV_X32 U_g21795 ( .A(I28314), .ZN(g21795) );
INV_X32 U_I28357 ( .A(g20497), .ZN(I28357) );
INV_X32 U_g21824 ( .A(I28357), .ZN(g21824) );
INV_X32 U_I28360 ( .A(g20163), .ZN(I28360) );
INV_X32 U_g21825 ( .A(I28360), .ZN(g21825) );
INV_X32 U_g21861 ( .A(g19657), .ZN(g21861) );
INV_X32 U_g21867 ( .A(g19705), .ZN(g21867) );
INV_X32 U_g21872 ( .A(g19749), .ZN(g21872) );
INV_X32 U_g21876 ( .A(g19792), .ZN(g21876) );
INV_X32 U_g21883 ( .A(g19890), .ZN(g21883) );
INV_X32 U_g21886 ( .A(g19915), .ZN(g21886) );
INV_X32 U_g21895 ( .A(g19945), .ZN(g21895) );
INV_X32 U_g21902 ( .A(g19978), .ZN(g21902) );
INV_X32 U_g21907 ( .A(g19972), .ZN(g21907) );
INV_X32 U_I28432 ( .A(g19335), .ZN(I28432) );
INV_X32 U_g21914 ( .A(I28432), .ZN(g21914) );
INV_X32 U_I28435 ( .A(g19358), .ZN(I28435) );
INV_X32 U_g21917 ( .A(I28435), .ZN(g21917) );
INV_X32 U_g21921 ( .A(g20002), .ZN(g21921) );
INV_X32 U_g21927 ( .A(g20045), .ZN(g21927) );
INV_X32 U_I28443 ( .A(g19358), .ZN(I28443) );
INV_X32 U_g21928 ( .A(I28443), .ZN(g21928) );
INV_X32 U_I28447 ( .A(g19369), .ZN(I28447) );
INV_X32 U_g21932 ( .A(I28447), .ZN(g21932) );
INV_X32 U_I28450 ( .A(g19390), .ZN(I28450) );
INV_X32 U_g21935 ( .A(I28450), .ZN(g21935) );
INV_X32 U_g21939 ( .A(g20040), .ZN(g21939) );
INV_X32 U_I28455 ( .A(g20943), .ZN(I28455) );
INV_X32 U_g21943 ( .A(I28455), .ZN(g21943) );
INV_X32 U_I28458 ( .A(g20971), .ZN(I28458) );
INV_X32 U_g21944 ( .A(I28458), .ZN(g21944) );
INV_X32 U_I28461 ( .A(g20998), .ZN(I28461) );
INV_X32 U_g21945 ( .A(I28461), .ZN(g21945) );
INV_X32 U_I28464 ( .A(g21024), .ZN(I28464) );
INV_X32 U_g21946 ( .A(I28464), .ZN(g21946) );
INV_X32 U_I28467 ( .A(g20942), .ZN(I28467) );
INV_X32 U_g21947 ( .A(I28467), .ZN(g21947) );
INV_X32 U_I28470 ( .A(g20984), .ZN(I28470) );
INV_X32 U_g21948 ( .A(I28470), .ZN(g21948) );
INV_X32 U_I28473 ( .A(g21030), .ZN(I28473) );
INV_X32 U_g21949 ( .A(I28473), .ZN(g21949) );
INV_X32 U_I28476 ( .A(g21064), .ZN(I28476) );
INV_X32 U_g21950 ( .A(I28476), .ZN(g21950) );
INV_X32 U_I28479 ( .A(g21795), .ZN(I28479) );
INV_X32 U_g21951 ( .A(I28479), .ZN(g21951) );
INV_X32 U_I28482 ( .A(g21376), .ZN(I28482) );
INV_X32 U_g21952 ( .A(I28482), .ZN(g21952) );
INV_X32 U_I28485 ( .A(g21426), .ZN(I28485) );
INV_X32 U_g21953 ( .A(I28485), .ZN(g21953) );
INV_X32 U_I28488 ( .A(g21495), .ZN(I28488) );
INV_X32 U_g21954 ( .A(I28488), .ZN(g21954) );
INV_X32 U_I28491 ( .A(g21327), .ZN(I28491) );
INV_X32 U_g21955 ( .A(I28491), .ZN(g21955) );
INV_X32 U_I28494 ( .A(g21358), .ZN(I28494) );
INV_X32 U_g21956 ( .A(I28494), .ZN(g21956) );
INV_X32 U_I28497 ( .A(g21399), .ZN(I28497) );
INV_X32 U_g21957 ( .A(I28497), .ZN(g21957) );
INV_X32 U_I28500 ( .A(g21457), .ZN(I28500) );
INV_X32 U_g21958 ( .A(I28500), .ZN(g21958) );
INV_X32 U_I28503 ( .A(g21528), .ZN(I28503) );
INV_X32 U_g21959 ( .A(I28503), .ZN(g21959) );
INV_X32 U_I28506 ( .A(g21377), .ZN(I28506) );
INV_X32 U_g21960 ( .A(I28506), .ZN(g21960) );
INV_X32 U_I28509 ( .A(g21427), .ZN(I28509) );
INV_X32 U_g21961 ( .A(I28509), .ZN(g21961) );
INV_X32 U_I28512 ( .A(g21496), .ZN(I28512) );
INV_X32 U_g21962 ( .A(I28512), .ZN(g21962) );
INV_X32 U_I28515 ( .A(g21557), .ZN(I28515) );
INV_X32 U_g21963 ( .A(I28515), .ZN(g21963) );
INV_X32 U_I28518 ( .A(g20985), .ZN(I28518) );
INV_X32 U_g21964 ( .A(I28518), .ZN(g21964) );
INV_X32 U_I28521 ( .A(g21824), .ZN(I28521) );
INV_X32 U_g21965 ( .A(I28521), .ZN(g21965) );
INV_X32 U_I28524 ( .A(g21359), .ZN(I28524) );
INV_X32 U_g21966 ( .A(I28524), .ZN(g21966) );
INV_X32 U_I28527 ( .A(g21407), .ZN(I28527) );
INV_X32 U_g21967 ( .A(I28527), .ZN(g21967) );
INV_X32 U_I28541 ( .A(g21467), .ZN(I28541) );
INV_X32 U_g21982 ( .A(I28541), .ZN(g21982) );
INV_X32 U_I28550 ( .A(g21432), .ZN(I28550) );
INV_X32 U_g21995 ( .A(I28550), .ZN(g21995) );
INV_X32 U_I28557 ( .A(g21407), .ZN(I28557) );
INV_X32 U_g22003 ( .A(I28557), .ZN(g22003) );
INV_X32 U_I28564 ( .A(g21385), .ZN(I28564) );
INV_X32 U_g22014 ( .A(I28564), .ZN(g22014) );
INV_X32 U_I28628 ( .A(g21842), .ZN(I28628) );
INV_X32 U_g22082 ( .A(I28628), .ZN(g22082) );
INV_X32 U_I28649 ( .A(g21843), .ZN(I28649) );
INV_X32 U_g22107 ( .A(I28649), .ZN(g22107) );
INV_X32 U_I28671 ( .A(g21845), .ZN(I28671) );
INV_X32 U_g22133 ( .A(I28671), .ZN(g22133) );
INV_X32 U_I28693 ( .A(g21847), .ZN(I28693) );
INV_X32 U_g22156 ( .A(I28693), .ZN(g22156) );
INV_X32 U_I28712 ( .A(g21851), .ZN(I28712) );
INV_X32 U_g22176 ( .A(I28712), .ZN(g22176) );
INV_X32 U_g22212 ( .A(g21914), .ZN(g22212) );
INV_X32 U_g22213 ( .A(g21917), .ZN(g22213) );
INV_X32 U_g22217 ( .A(g21928), .ZN(g22217) );
INV_X32 U_I28781 ( .A(g21331), .ZN(I28781) );
INV_X32 U_g22219 ( .A(I28781), .ZN(g22219) );
INV_X32 U_g22221 ( .A(g21932), .ZN(g22221) );
INV_X32 U_g22222 ( .A(g21935), .ZN(g22222) );
INV_X32 U_I28789 ( .A(g21878), .ZN(I28789) );
INV_X32 U_g22225 ( .A(I28789), .ZN(g22225) );
INV_X32 U_I28792 ( .A(g21880), .ZN(I28792) );
INV_X32 U_g22226 ( .A(I28792), .ZN(g22226) );
INV_X32 U_g22230 ( .A(g20634), .ZN(g22230) );
INV_X32 U_I28800 ( .A(g21316), .ZN(I28800) );
INV_X32 U_g22232 ( .A(I28800), .ZN(g22232) );
INV_X32 U_g22233 ( .A(g20637), .ZN(g22233) );
INV_X32 U_g22236 ( .A(g20641), .ZN(g22236) );
INV_X32 U_g22237 ( .A(g20644), .ZN(g22237) );
INV_X32 U_g22239 ( .A(g20649), .ZN(g22239) );
INV_X32 U_g22240 ( .A(g20652), .ZN(g22240) );
INV_X32 U_g22241 ( .A(g20655), .ZN(g22241) );
INV_X32 U_I28813 ( .A(g21502), .ZN(I28813) );
INV_X32 U_g22243 ( .A(I28813), .ZN(g22243) );
INV_X32 U_g22246 ( .A(g20659), .ZN(g22246) );
INV_X32 U_g22248 ( .A(g20662), .ZN(g22248) );
INV_X32 U_g22251 ( .A(g20666), .ZN(g22251) );
INV_X32 U_g22252 ( .A(g20669), .ZN(g22252) );
INV_X32 U_I28825 ( .A(g21882), .ZN(I28825) );
INV_X32 U_g22253 ( .A(I28825), .ZN(g22253) );
INV_X32 U_g22256 ( .A(g20673), .ZN(g22256) );
INV_X32 U_g22257 ( .A(g20676), .ZN(g22257) );
INV_X32 U_g22258 ( .A(g20679), .ZN(g22258) );
INV_X32 U_I28833 ( .A(g21470), .ZN(I28833) );
INV_X32 U_g22259 ( .A(I28833), .ZN(g22259) );
INV_X32 U_g22260 ( .A(g20684), .ZN(g22260) );
INV_X32 U_g22261 ( .A(g20687), .ZN(g22261) );
INV_X32 U_g22262 ( .A(g20690), .ZN(g22262) );
INV_X32 U_g22266 ( .A(g20694), .ZN(g22266) );
INV_X32 U_g22268 ( .A(g20697), .ZN(g22268) );
INV_X32 U_g22271 ( .A(g20704), .ZN(g22271) );
INV_X32 U_g22274 ( .A(g20708), .ZN(g22274) );
INV_X32 U_g22275 ( .A(g20711), .ZN(g22275) );
INV_X32 U_g22276 ( .A(g20714), .ZN(g22276) );
INV_X32 U_g22277 ( .A(g20719), .ZN(g22277) );
INV_X32 U_g22278 ( .A(g20722), .ZN(g22278) );
INV_X32 U_g22279 ( .A(g20725), .ZN(g22279) );
INV_X32 U_g22283 ( .A(g20729), .ZN(g22283) );
INV_X32 U_g22286 ( .A(g20732), .ZN(g22286) );
INV_X32 U_g22287 ( .A(g20735), .ZN(g22287) );
INV_X32 U_g22290 ( .A(g20739), .ZN(g22290) );
INV_X32 U_g22293 ( .A(g20743), .ZN(g22293) );
INV_X32 U_g22294 ( .A(g20746), .ZN(g22294) );
INV_X32 U_g22295 ( .A(g20749), .ZN(g22295) );
INV_X32 U_g22296 ( .A(g20754), .ZN(g22296) );
INV_X32 U_g22297 ( .A(g20757), .ZN(g22297) );
INV_X32 U_g22298 ( .A(g20760), .ZN(g22298) );
INV_X32 U_I28876 ( .A(g21238), .ZN(I28876) );
INV_X32 U_g22300 ( .A(I28876), .ZN(g22300) );
INV_X32 U_g22303 ( .A(g20763), .ZN(g22303) );
INV_X32 U_g22304 ( .A(g20766), .ZN(g22304) );
INV_X32 U_g22306 ( .A(g20769), .ZN(g22306) );
INV_X32 U_g22307 ( .A(g20772), .ZN(g22307) );
INV_X32 U_g22310 ( .A(g20776), .ZN(g22310) );
INV_X32 U_g22313 ( .A(g20780), .ZN(g22313) );
INV_X32 U_g22314 ( .A(g20783), .ZN(g22314) );
INV_X32 U_g22315 ( .A(g20786), .ZN(g22315) );
INV_X32 U_g22316 ( .A(g21149), .ZN(g22316) );
INV_X32 U_g22318 ( .A(g20790), .ZN(g22318) );
INV_X32 U_g22319 ( .A(g21228), .ZN(g22319) );
INV_X32 U_I28896 ( .A(g21246), .ZN(I28896) );
INV_X32 U_g22328 ( .A(I28896), .ZN(g22328) );
INV_X32 U_g22331 ( .A(g20793), .ZN(g22331) );
INV_X32 U_g22332 ( .A(g20796), .ZN(g22332) );
INV_X32 U_g22334 ( .A(g20799), .ZN(g22334) );
INV_X32 U_g22335 ( .A(g20802), .ZN(g22335) );
INV_X32 U_g22338 ( .A(g20806), .ZN(g22338) );
INV_X32 U_g22341 ( .A(g21169), .ZN(g22341) );
INV_X32 U_g22343 ( .A(g20810), .ZN(g22343) );
INV_X32 U_g22344 ( .A(g21233), .ZN(g22344) );
INV_X32 U_I28913 ( .A(g21255), .ZN(I28913) );
INV_X32 U_g22353 ( .A(I28913), .ZN(g22353) );
INV_X32 U_g22356 ( .A(g20813), .ZN(g22356) );
INV_X32 U_g22357 ( .A(g20816), .ZN(g22357) );
INV_X32 U_g22359 ( .A(g20819), .ZN(g22359) );
INV_X32 U_g22360 ( .A(g20822), .ZN(g22360) );
INV_X32 U_g22364 ( .A(g21189), .ZN(g22364) );
INV_X32 U_g22366 ( .A(g20827), .ZN(g22366) );
INV_X32 U_g22367 ( .A(g21242), .ZN(g22367) );
INV_X32 U_I28928 ( .A(g21263), .ZN(I28928) );
INV_X32 U_g22376 ( .A(I28928), .ZN(g22376) );
INV_X32 U_g22379 ( .A(g20830), .ZN(g22379) );
INV_X32 U_g22380 ( .A(g20833), .ZN(g22380) );
INV_X32 U_g22384 ( .A(g21204), .ZN(g22384) );
INV_X32 U_g22386 ( .A(g20837), .ZN(g22386) );
INV_X32 U_g22387 ( .A(g21250), .ZN(g22387) );
INV_X32 U_g22401 ( .A(g21533), .ZN(g22401) );
INV_X32 U_g22402 ( .A(g21569), .ZN(g22402) );
INV_X32 U_g22403 ( .A(g21602), .ZN(g22403) );
INV_X32 U_g22404 ( .A(g21631), .ZN(g22404) );
INV_X32 U_I28949 ( .A(g21685), .ZN(I28949) );
INV_X32 U_g22405 ( .A(I28949), .ZN(g22405) );
INV_X32 U_g22408 ( .A(g20986), .ZN(g22408) );
INV_X32 U_I28953 ( .A(g21659), .ZN(I28953) );
INV_X32 U_g22409 ( .A(I28953), .ZN(g22409) );
INV_X32 U_I28956 ( .A(g21714), .ZN(I28956) );
INV_X32 U_g22412 ( .A(I28956), .ZN(g22412) );
INV_X32 U_I28959 ( .A(g21636), .ZN(I28959) );
INV_X32 U_g22415 ( .A(I28959), .ZN(g22415) );
INV_X32 U_I28962 ( .A(g21721), .ZN(I28962) );
INV_X32 U_g22418 ( .A(I28962), .ZN(g22418) );
INV_X32 U_g22421 ( .A(g21012), .ZN(g22421) );
INV_X32 U_I28966 ( .A(g20633), .ZN(I28966) );
INV_X32 U_g22422 ( .A(I28966), .ZN(g22422) );
INV_X32 U_I28969 ( .A(g21686), .ZN(I28969) );
INV_X32 U_g22425 ( .A(I28969), .ZN(g22425) );
INV_X32 U_I28972 ( .A(g21736), .ZN(I28972) );
INV_X32 U_g22428 ( .A(I28972), .ZN(g22428) );
INV_X32 U_I28975 ( .A(g21688), .ZN(I28975) );
INV_X32 U_g22431 ( .A(I28975), .ZN(g22431) );
INV_X32 U_I28978 ( .A(g21740), .ZN(I28978) );
INV_X32 U_g22434 ( .A(I28978), .ZN(g22434) );
INV_X32 U_I28981 ( .A(g21667), .ZN(I28981) );
INV_X32 U_g22437 ( .A(I28981), .ZN(g22437) );
INV_X32 U_I28984 ( .A(g21747), .ZN(I28984) );
INV_X32 U_g22440 ( .A(I28984), .ZN(g22440) );
INV_X32 U_g22443 ( .A(g21036), .ZN(g22443) );
INV_X32 U_I28988 ( .A(g20874), .ZN(I28988) );
INV_X32 U_g22444 ( .A(I28988), .ZN(g22444) );
INV_X32 U_I28991 ( .A(g20648), .ZN(I28991) );
INV_X32 U_g22445 ( .A(I28991), .ZN(g22445) );
INV_X32 U_I28994 ( .A(g21715), .ZN(I28994) );
INV_X32 U_g22448 ( .A(I28994), .ZN(g22448) );
INV_X32 U_I28997 ( .A(g21759), .ZN(I28997) );
INV_X32 U_g22451 ( .A(I28997), .ZN(g22451) );
INV_X32 U_I29001 ( .A(g20658), .ZN(I29001) );
INV_X32 U_g22455 ( .A(I29001), .ZN(g22455) );
INV_X32 U_I29004 ( .A(g21722), .ZN(I29004) );
INV_X32 U_g22458 ( .A(I29004), .ZN(g22458) );
INV_X32 U_I29007 ( .A(g21760), .ZN(I29007) );
INV_X32 U_g22461 ( .A(I29007), .ZN(g22461) );
INV_X32 U_I29010 ( .A(g21724), .ZN(I29010) );
INV_X32 U_g22464 ( .A(I29010), .ZN(g22464) );
INV_X32 U_I29013 ( .A(g21764), .ZN(I29013) );
INV_X32 U_g22467 ( .A(I29013), .ZN(g22467) );
INV_X32 U_I29016 ( .A(g21696), .ZN(I29016) );
INV_X32 U_g22470 ( .A(I29016), .ZN(g22470) );
INV_X32 U_I29019 ( .A(g21771), .ZN(I29019) );
INV_X32 U_g22473 ( .A(I29019), .ZN(g22473) );
INV_X32 U_g22476 ( .A(g21057), .ZN(g22476) );
INV_X32 U_I29023 ( .A(g20672), .ZN(I29023) );
INV_X32 U_g22477 ( .A(I29023), .ZN(g22477) );
INV_X32 U_I29026 ( .A(g21737), .ZN(I29026) );
INV_X32 U_g22480 ( .A(I29026), .ZN(g22480) );
INV_X32 U_I29030 ( .A(g20683), .ZN(I29030) );
INV_X32 U_g22484 ( .A(I29030), .ZN(g22484) );
INV_X32 U_I29033 ( .A(g21741), .ZN(I29033) );
INV_X32 U_g22487 ( .A(I29033), .ZN(g22487) );
INV_X32 U_I29036 ( .A(g21775), .ZN(I29036) );
INV_X32 U_g22490 ( .A(I29036), .ZN(g22490) );
INV_X32 U_I29040 ( .A(g20693), .ZN(I29040) );
INV_X32 U_g22494 ( .A(I29040), .ZN(g22494) );
INV_X32 U_I29043 ( .A(g21748), .ZN(I29043) );
INV_X32 U_g22497 ( .A(I29043), .ZN(g22497) );
INV_X32 U_I29046 ( .A(g21776), .ZN(I29046) );
INV_X32 U_g22500 ( .A(I29046), .ZN(g22500) );
INV_X32 U_I29049 ( .A(g21750), .ZN(I29049) );
INV_X32 U_g22503 ( .A(I29049), .ZN(g22503) );
INV_X32 U_I29052 ( .A(g21780), .ZN(I29052) );
INV_X32 U_g22506 ( .A(I29052), .ZN(g22506) );
INV_X32 U_I29055 ( .A(g21732), .ZN(I29055) );
INV_X32 U_g22509 ( .A(I29055), .ZN(g22509) );
INV_X32 U_I29058 ( .A(g20703), .ZN(I29058) );
INV_X32 U_g22512 ( .A(I29058), .ZN(g22512) );
INV_X32 U_I29064 ( .A(g20875), .ZN(I29064) );
INV_X32 U_g22518 ( .A(I29064), .ZN(g22518) );
INV_X32 U_I29067 ( .A(g20876), .ZN(I29067) );
INV_X32 U_g22519 ( .A(I29067), .ZN(g22519) );
INV_X32 U_I29070 ( .A(g20707), .ZN(I29070) );
INV_X32 U_g22520 ( .A(I29070), .ZN(g22520) );
INV_X32 U_I29073 ( .A(g21761), .ZN(I29073) );
INV_X32 U_g22523 ( .A(I29073), .ZN(g22523) );
INV_X32 U_I29077 ( .A(g20718), .ZN(I29077) );
INV_X32 U_g22527 ( .A(I29077), .ZN(g22527) );
INV_X32 U_I29080 ( .A(g21765), .ZN(I29080) );
INV_X32 U_g22530 ( .A(I29080), .ZN(g22530) );
INV_X32 U_I29083 ( .A(g21790), .ZN(I29083) );
INV_X32 U_g22533 ( .A(I29083), .ZN(g22533) );
INV_X32 U_I29087 ( .A(g20728), .ZN(I29087) );
INV_X32 U_g22537 ( .A(I29087), .ZN(g22537) );
INV_X32 U_I29090 ( .A(g21772), .ZN(I29090) );
INV_X32 U_g22540 ( .A(I29090), .ZN(g22540) );
INV_X32 U_I29093 ( .A(g21791), .ZN(I29093) );
INV_X32 U_g22543 ( .A(I29093), .ZN(g22543) );
INV_X32 U_g22547 ( .A(g21087), .ZN(g22547) );
INV_X32 U_I29098 ( .A(g20879), .ZN(I29098) );
INV_X32 U_g22548 ( .A(I29098), .ZN(g22548) );
INV_X32 U_I29101 ( .A(g20880), .ZN(I29101) );
INV_X32 U_g22549 ( .A(I29101), .ZN(g22549) );
INV_X32 U_I29104 ( .A(g20881), .ZN(I29104) );
INV_X32 U_g22550 ( .A(I29104), .ZN(g22550) );
INV_X32 U_I29107 ( .A(g21435), .ZN(I29107) );
INV_X32 U_g22551 ( .A(I29107), .ZN(g22551) );
INV_X32 U_I29110 ( .A(g20738), .ZN(I29110) );
INV_X32 U_g22552 ( .A(I29110), .ZN(g22552) );
INV_X32 U_I29116 ( .A(g20882), .ZN(I29116) );
INV_X32 U_g22558 ( .A(I29116), .ZN(g22558) );
INV_X32 U_I29119 ( .A(g20883), .ZN(I29119) );
INV_X32 U_g22559 ( .A(I29119), .ZN(g22559) );
INV_X32 U_I29122 ( .A(g20742), .ZN(I29122) );
INV_X32 U_g22560 ( .A(I29122), .ZN(g22560) );
INV_X32 U_I29125 ( .A(g21777), .ZN(I29125) );
INV_X32 U_g22563 ( .A(I29125), .ZN(g22563) );
INV_X32 U_I29129 ( .A(g20753), .ZN(I29129) );
INV_X32 U_g22567 ( .A(I29129), .ZN(g22567) );
INV_X32 U_I29132 ( .A(g21781), .ZN(I29132) );
INV_X32 U_g22570 ( .A(I29132), .ZN(g22570) );
INV_X32 U_I29135 ( .A(g21804), .ZN(I29135) );
INV_X32 U_g22573 ( .A(I29135), .ZN(g22573) );
INV_X32 U_I29142 ( .A(g20682), .ZN(I29142) );
INV_X32 U_g22582 ( .A(I29142), .ZN(g22582) );
INV_X32 U_I29145 ( .A(g20891), .ZN(I29145) );
INV_X32 U_g22583 ( .A(I29145), .ZN(g22583) );
INV_X32 U_I29148 ( .A(g20892), .ZN(I29148) );
INV_X32 U_g22584 ( .A(I29148), .ZN(g22584) );
INV_X32 U_I29151 ( .A(g20893), .ZN(I29151) );
INV_X32 U_g22585 ( .A(I29151), .ZN(g22585) );
INV_X32 U_I29154 ( .A(g20894), .ZN(I29154) );
INV_X32 U_g22586 ( .A(I29154), .ZN(g22586) );
INV_X32 U_g22588 ( .A(g21099), .ZN(g22588) );
INV_X32 U_I29159 ( .A(g20896), .ZN(I29159) );
INV_X32 U_g22589 ( .A(I29159), .ZN(g22589) );
INV_X32 U_I29162 ( .A(g20897), .ZN(I29162) );
INV_X32 U_g22590 ( .A(I29162), .ZN(g22590) );
INV_X32 U_I29165 ( .A(g20898), .ZN(I29165) );
INV_X32 U_g22591 ( .A(I29165), .ZN(g22591) );
INV_X32 U_I29168 ( .A(g20775), .ZN(I29168) );
INV_X32 U_g22592 ( .A(I29168), .ZN(g22592) );
INV_X32 U_I29174 ( .A(g20899), .ZN(I29174) );
INV_X32 U_g22598 ( .A(I29174), .ZN(g22598) );
INV_X32 U_I29177 ( .A(g20900), .ZN(I29177) );
INV_X32 U_g22599 ( .A(I29177), .ZN(g22599) );
INV_X32 U_I29180 ( .A(g20779), .ZN(I29180) );
INV_X32 U_g22600 ( .A(I29180), .ZN(g22600) );
INV_X32 U_I29183 ( .A(g21792), .ZN(I29183) );
INV_X32 U_g22603 ( .A(I29183), .ZN(g22603) );
INV_X32 U_g22609 ( .A(g21108), .ZN(g22609) );
INV_X32 U_I29191 ( .A(g20901), .ZN(I29191) );
INV_X32 U_g22611 ( .A(I29191), .ZN(g22611) );
INV_X32 U_I29194 ( .A(g20902), .ZN(I29194) );
INV_X32 U_g22612 ( .A(I29194), .ZN(g22612) );
INV_X32 U_I29197 ( .A(g20903), .ZN(I29197) );
INV_X32 U_g22613 ( .A(I29197), .ZN(g22613) );
INV_X32 U_I29203 ( .A(g20717), .ZN(I29203) );
INV_X32 U_g22619 ( .A(I29203), .ZN(g22619) );
INV_X32 U_I29206 ( .A(g20910), .ZN(I29206) );
INV_X32 U_g22620 ( .A(I29206), .ZN(g22620) );
INV_X32 U_I29209 ( .A(g20911), .ZN(I29209) );
INV_X32 U_g22621 ( .A(I29209), .ZN(g22621) );
INV_X32 U_I29212 ( .A(g20912), .ZN(I29212) );
INV_X32 U_g22622 ( .A(I29212), .ZN(g22622) );
INV_X32 U_I29215 ( .A(g20913), .ZN(I29215) );
INV_X32 U_g22623 ( .A(I29215), .ZN(g22623) );
INV_X32 U_g22625 ( .A(g21113), .ZN(g22625) );
INV_X32 U_I29220 ( .A(g20915), .ZN(I29220) );
INV_X32 U_g22626 ( .A(I29220), .ZN(g22626) );
INV_X32 U_I29223 ( .A(g20916), .ZN(I29223) );
INV_X32 U_g22627 ( .A(I29223), .ZN(g22627) );
INV_X32 U_I29226 ( .A(g20917), .ZN(I29226) );
INV_X32 U_g22628 ( .A(I29226), .ZN(g22628) );
INV_X32 U_I29229 ( .A(g20805), .ZN(I29229) );
INV_X32 U_g22629 ( .A(I29229), .ZN(g22629) );
INV_X32 U_I29235 ( .A(g20918), .ZN(I29235) );
INV_X32 U_g22635 ( .A(I29235), .ZN(g22635) );
INV_X32 U_I29238 ( .A(g20919), .ZN(I29238) );
INV_X32 U_g22636 ( .A(I29238), .ZN(g22636) );
INV_X32 U_I29243 ( .A(g20921), .ZN(I29243) );
INV_X32 U_g22639 ( .A(I29243), .ZN(g22639) );
INV_X32 U_I29246 ( .A(g20922), .ZN(I29246) );
INV_X32 U_g22640 ( .A(I29246), .ZN(g22640) );
INV_X32 U_I29249 ( .A(g20923), .ZN(I29249) );
INV_X32 U_g22641 ( .A(I29249), .ZN(g22641) );
INV_X32 U_I29252 ( .A(g20924), .ZN(I29252) );
INV_X32 U_g22642 ( .A(I29252), .ZN(g22642) );
INV_X32 U_g22645 ( .A(g21125), .ZN(g22645) );
INV_X32 U_I29259 ( .A(g20925), .ZN(I29259) );
INV_X32 U_g22647 ( .A(I29259), .ZN(g22647) );
INV_X32 U_I29262 ( .A(g20926), .ZN(I29262) );
INV_X32 U_g22648 ( .A(I29262), .ZN(g22648) );
INV_X32 U_I29265 ( .A(g20927), .ZN(I29265) );
INV_X32 U_g22649 ( .A(I29265), .ZN(g22649) );
INV_X32 U_I29271 ( .A(g20752), .ZN(I29271) );
INV_X32 U_g22655 ( .A(I29271), .ZN(g22655) );
INV_X32 U_I29274 ( .A(g20934), .ZN(I29274) );
INV_X32 U_g22656 ( .A(I29274), .ZN(g22656) );
INV_X32 U_I29277 ( .A(g20935), .ZN(I29277) );
INV_X32 U_g22657 ( .A(I29277), .ZN(g22657) );
INV_X32 U_I29280 ( .A(g20936), .ZN(I29280) );
INV_X32 U_g22658 ( .A(I29280), .ZN(g22658) );
INV_X32 U_I29283 ( .A(g20937), .ZN(I29283) );
INV_X32 U_g22659 ( .A(I29283), .ZN(g22659) );
INV_X32 U_g22661 ( .A(g21130), .ZN(g22661) );
INV_X32 U_I29288 ( .A(g20939), .ZN(I29288) );
INV_X32 U_g22662 ( .A(I29288), .ZN(g22662) );
INV_X32 U_I29291 ( .A(g20940), .ZN(I29291) );
INV_X32 U_g22663 ( .A(I29291), .ZN(g22663) );
INV_X32 U_I29294 ( .A(g20941), .ZN(I29294) );
INV_X32 U_g22664 ( .A(I29294), .ZN(g22664) );
INV_X32 U_I29301 ( .A(g20944), .ZN(I29301) );
INV_X32 U_g22669 ( .A(I29301), .ZN(g22669) );
INV_X32 U_I29304 ( .A(g20945), .ZN(I29304) );
INV_X32 U_g22670 ( .A(I29304), .ZN(g22670) );
INV_X32 U_I29307 ( .A(g20946), .ZN(I29307) );
INV_X32 U_g22671 ( .A(I29307), .ZN(g22671) );
INV_X32 U_I29310 ( .A(g20947), .ZN(I29310) );
INV_X32 U_g22672 ( .A(I29310), .ZN(g22672) );
INV_X32 U_I29313 ( .A(g20948), .ZN(I29313) );
INV_X32 U_g22673 ( .A(I29313), .ZN(g22673) );
INV_X32 U_I29317 ( .A(g20949), .ZN(I29317) );
INV_X32 U_g22675 ( .A(I29317), .ZN(g22675) );
INV_X32 U_I29320 ( .A(g20950), .ZN(I29320) );
INV_X32 U_g22676 ( .A(I29320), .ZN(g22676) );
INV_X32 U_I29323 ( .A(g20951), .ZN(I29323) );
INV_X32 U_g22677 ( .A(I29323), .ZN(g22677) );
INV_X32 U_I29326 ( .A(g20952), .ZN(I29326) );
INV_X32 U_g22678 ( .A(I29326), .ZN(g22678) );
INV_X32 U_g22681 ( .A(g21144), .ZN(g22681) );
INV_X32 U_I29333 ( .A(g20953), .ZN(I29333) );
INV_X32 U_g22683 ( .A(I29333), .ZN(g22683) );
INV_X32 U_I29336 ( .A(g20954), .ZN(I29336) );
INV_X32 U_g22684 ( .A(I29336), .ZN(g22684) );
INV_X32 U_I29339 ( .A(g20955), .ZN(I29339) );
INV_X32 U_g22685 ( .A(I29339), .ZN(g22685) );
INV_X32 U_I29345 ( .A(g20789), .ZN(I29345) );
INV_X32 U_g22691 ( .A(I29345), .ZN(g22691) );
INV_X32 U_I29348 ( .A(g20962), .ZN(I29348) );
INV_X32 U_g22692 ( .A(I29348), .ZN(g22692) );
INV_X32 U_I29351 ( .A(g20963), .ZN(I29351) );
INV_X32 U_g22693 ( .A(I29351), .ZN(g22693) );
INV_X32 U_I29354 ( .A(g20964), .ZN(I29354) );
INV_X32 U_g22694 ( .A(I29354), .ZN(g22694) );
INV_X32 U_I29357 ( .A(g20965), .ZN(I29357) );
INV_X32 U_g22695 ( .A(I29357), .ZN(g22695) );
INV_X32 U_I29360 ( .A(g21796), .ZN(I29360) );
INV_X32 U_g22696 ( .A(I29360), .ZN(g22696) );
INV_X32 U_I29366 ( .A(g20966), .ZN(I29366) );
INV_X32 U_g22702 ( .A(I29366), .ZN(g22702) );
INV_X32 U_I29369 ( .A(g20967), .ZN(I29369) );
INV_X32 U_g22703 ( .A(I29369), .ZN(g22703) );
INV_X32 U_I29372 ( .A(g20968), .ZN(I29372) );
INV_X32 U_g22704 ( .A(I29372), .ZN(g22704) );
INV_X32 U_I29375 ( .A(g20969), .ZN(I29375) );
INV_X32 U_g22705 ( .A(I29375), .ZN(g22705) );
INV_X32 U_I29378 ( .A(g20970), .ZN(I29378) );
INV_X32 U_g22706 ( .A(I29378), .ZN(g22706) );
INV_X32 U_I29383 ( .A(g20972), .ZN(I29383) );
INV_X32 U_g22709 ( .A(I29383), .ZN(g22709) );
INV_X32 U_I29386 ( .A(g20973), .ZN(I29386) );
INV_X32 U_g22710 ( .A(I29386), .ZN(g22710) );
INV_X32 U_I29389 ( .A(g20974), .ZN(I29389) );
INV_X32 U_g22711 ( .A(I29389), .ZN(g22711) );
INV_X32 U_I29392 ( .A(g20975), .ZN(I29392) );
INV_X32 U_g22712 ( .A(I29392), .ZN(g22712) );
INV_X32 U_I29395 ( .A(g20976), .ZN(I29395) );
INV_X32 U_g22713 ( .A(I29395), .ZN(g22713) );
INV_X32 U_I29399 ( .A(g20977), .ZN(I29399) );
INV_X32 U_g22715 ( .A(I29399), .ZN(g22715) );
INV_X32 U_I29402 ( .A(g20978), .ZN(I29402) );
INV_X32 U_g22716 ( .A(I29402), .ZN(g22716) );
INV_X32 U_I29405 ( .A(g20979), .ZN(I29405) );
INV_X32 U_g22717 ( .A(I29405), .ZN(g22717) );
INV_X32 U_I29408 ( .A(g20980), .ZN(I29408) );
INV_X32 U_g22718 ( .A(I29408), .ZN(g22718) );
INV_X32 U_g22721 ( .A(g21164), .ZN(g22721) );
INV_X32 U_I29415 ( .A(g20981), .ZN(I29415) );
INV_X32 U_g22723 ( .A(I29415), .ZN(g22723) );
INV_X32 U_I29418 ( .A(g20982), .ZN(I29418) );
INV_X32 U_g22724 ( .A(I29418), .ZN(g22724) );
INV_X32 U_I29421 ( .A(g20983), .ZN(I29421) );
INV_X32 U_g22725 ( .A(I29421), .ZN(g22725) );
INV_X32 U_I29426 ( .A(g20989), .ZN(I29426) );
INV_X32 U_g22728 ( .A(I29426), .ZN(g22728) );
INV_X32 U_I29429 ( .A(g20990), .ZN(I29429) );
INV_X32 U_g22729 ( .A(I29429), .ZN(g22729) );
INV_X32 U_I29432 ( .A(g20991), .ZN(I29432) );
INV_X32 U_g22730 ( .A(I29432), .ZN(g22730) );
INV_X32 U_I29435 ( .A(g20992), .ZN(I29435) );
INV_X32 U_g22731 ( .A(I29435), .ZN(g22731) );
INV_X32 U_I29439 ( .A(g20993), .ZN(I29439) );
INV_X32 U_g22733 ( .A(I29439), .ZN(g22733) );
INV_X32 U_I29442 ( .A(g20994), .ZN(I29442) );
INV_X32 U_g22734 ( .A(I29442), .ZN(g22734) );
INV_X32 U_I29445 ( .A(g20995), .ZN(I29445) );
INV_X32 U_g22735 ( .A(I29445), .ZN(g22735) );
INV_X32 U_I29448 ( .A(g20996), .ZN(I29448) );
INV_X32 U_g22736 ( .A(I29448), .ZN(g22736) );
INV_X32 U_I29451 ( .A(g20997), .ZN(I29451) );
INV_X32 U_g22737 ( .A(I29451), .ZN(g22737) );
INV_X32 U_I29456 ( .A(g20999), .ZN(I29456) );
INV_X32 U_g22740 ( .A(I29456), .ZN(g22740) );
INV_X32 U_I29459 ( .A(g21000), .ZN(I29459) );
INV_X32 U_g22741 ( .A(I29459), .ZN(g22741) );
INV_X32 U_I29462 ( .A(g21001), .ZN(I29462) );
INV_X32 U_g22742 ( .A(I29462), .ZN(g22742) );
INV_X32 U_I29465 ( .A(g21002), .ZN(I29465) );
INV_X32 U_g22743 ( .A(I29465), .ZN(g22743) );
INV_X32 U_I29468 ( .A(g21003), .ZN(I29468) );
INV_X32 U_g22744 ( .A(I29468), .ZN(g22744) );
INV_X32 U_I29472 ( .A(g21004), .ZN(I29472) );
INV_X32 U_g22746 ( .A(I29472), .ZN(g22746) );
INV_X32 U_I29475 ( .A(g21005), .ZN(I29475) );
INV_X32 U_g22747 ( .A(I29475), .ZN(g22747) );
INV_X32 U_I29478 ( .A(g21006), .ZN(I29478) );
INV_X32 U_g22748 ( .A(I29478), .ZN(g22748) );
INV_X32 U_I29481 ( .A(g21007), .ZN(I29481) );
INV_X32 U_g22749 ( .A(I29481), .ZN(g22749) );
INV_X32 U_I29484 ( .A(g21903), .ZN(I29484) );
INV_X32 U_g22750 ( .A(I29484), .ZN(g22750) );
INV_X32 U_g22753 ( .A(g21184), .ZN(g22753) );
INV_X32 U_I29490 ( .A(g21009), .ZN(I29490) );
INV_X32 U_g22756 ( .A(I29490), .ZN(g22756) );
INV_X32 U_I29493 ( .A(g21010), .ZN(I29493) );
INV_X32 U_g22757 ( .A(I29493), .ZN(g22757) );
INV_X32 U_I29496 ( .A(g21011), .ZN(I29496) );
INV_X32 U_g22758 ( .A(I29496), .ZN(g22758) );
INV_X32 U_I29500 ( .A(g21015), .ZN(I29500) );
INV_X32 U_g22760 ( .A(I29500), .ZN(g22760) );
INV_X32 U_I29503 ( .A(g21016), .ZN(I29503) );
INV_X32 U_g22761 ( .A(I29503), .ZN(g22761) );
INV_X32 U_I29506 ( .A(g21017), .ZN(I29506) );
INV_X32 U_g22762 ( .A(I29506), .ZN(g22762) );
INV_X32 U_I29509 ( .A(g21018), .ZN(I29509) );
INV_X32 U_g22763 ( .A(I29509), .ZN(g22763) );
INV_X32 U_I29513 ( .A(g21019), .ZN(I29513) );
INV_X32 U_g22765 ( .A(I29513), .ZN(g22765) );
INV_X32 U_I29516 ( .A(g21020), .ZN(I29516) );
INV_X32 U_g22766 ( .A(I29516), .ZN(g22766) );
INV_X32 U_I29519 ( .A(g21021), .ZN(I29519) );
INV_X32 U_g22767 ( .A(I29519), .ZN(g22767) );
INV_X32 U_I29522 ( .A(g21022), .ZN(I29522) );
INV_X32 U_g22768 ( .A(I29522), .ZN(g22768) );
INV_X32 U_I29525 ( .A(g21023), .ZN(I29525) );
INV_X32 U_g22769 ( .A(I29525), .ZN(g22769) );
INV_X32 U_I29530 ( .A(g21025), .ZN(I29530) );
INV_X32 U_g22772 ( .A(I29530), .ZN(g22772) );
INV_X32 U_I29533 ( .A(g21026), .ZN(I29533) );
INV_X32 U_g22773 ( .A(I29533), .ZN(g22773) );
INV_X32 U_I29536 ( .A(g21027), .ZN(I29536) );
INV_X32 U_g22774 ( .A(I29536), .ZN(g22774) );
INV_X32 U_I29539 ( .A(g21028), .ZN(I29539) );
INV_X32 U_g22775 ( .A(I29539), .ZN(g22775) );
INV_X32 U_I29542 ( .A(g21029), .ZN(I29542) );
INV_X32 U_g22776 ( .A(I29542), .ZN(g22776) );
INV_X32 U_g22777 ( .A(g21796), .ZN(g22777) );
INV_X32 U_I29547 ( .A(g21031), .ZN(I29547) );
INV_X32 U_g22785 ( .A(I29547), .ZN(g22785) );
INV_X32 U_I29550 ( .A(g21032), .ZN(I29550) );
INV_X32 U_g22786 ( .A(I29550), .ZN(g22786) );
INV_X32 U_g22787 ( .A(g21199), .ZN(g22787) );
INV_X32 U_I29556 ( .A(g21033), .ZN(I29556) );
INV_X32 U_g22790 ( .A(I29556), .ZN(g22790) );
INV_X32 U_I29559 ( .A(g21034), .ZN(I29559) );
INV_X32 U_g22791 ( .A(I29559), .ZN(g22791) );
INV_X32 U_I29562 ( .A(g21035), .ZN(I29562) );
INV_X32 U_g22792 ( .A(I29562), .ZN(g22792) );
INV_X32 U_I29566 ( .A(g21039), .ZN(I29566) );
INV_X32 U_g22794 ( .A(I29566), .ZN(g22794) );
INV_X32 U_I29569 ( .A(g21040), .ZN(I29569) );
INV_X32 U_g22795 ( .A(I29569), .ZN(g22795) );
INV_X32 U_I29572 ( .A(g21041), .ZN(I29572) );
INV_X32 U_g22796 ( .A(I29572), .ZN(g22796) );
INV_X32 U_I29575 ( .A(g21042), .ZN(I29575) );
INV_X32 U_g22797 ( .A(I29575), .ZN(g22797) );
INV_X32 U_I29579 ( .A(g21043), .ZN(I29579) );
INV_X32 U_g22799 ( .A(I29579), .ZN(g22799) );
INV_X32 U_I29582 ( .A(g21044), .ZN(I29582) );
INV_X32 U_g22800 ( .A(I29582), .ZN(g22800) );
INV_X32 U_I29585 ( .A(g21045), .ZN(I29585) );
INV_X32 U_g22801 ( .A(I29585), .ZN(g22801) );
INV_X32 U_I29588 ( .A(g21046), .ZN(I29588) );
INV_X32 U_g22802 ( .A(I29588), .ZN(g22802) );
INV_X32 U_I29591 ( .A(g21047), .ZN(I29591) );
INV_X32 U_g22803 ( .A(I29591), .ZN(g22803) );
INV_X32 U_g22805 ( .A(g21894), .ZN(g22805) );
INV_X32 U_g22806 ( .A(g21615), .ZN(g22806) );
INV_X32 U_I29600 ( .A(g21720), .ZN(I29600) );
INV_X32 U_g22812 ( .A(I29600), .ZN(g22812) );
INV_X32 U_I29603 ( .A(g21051), .ZN(I29603) );
INV_X32 U_g22824 ( .A(I29603), .ZN(g22824) );
INV_X32 U_I29606 ( .A(g21364), .ZN(I29606) );
INV_X32 U_g22825 ( .A(I29606), .ZN(g22825) );
INV_X32 U_I29610 ( .A(g21052), .ZN(I29610) );
INV_X32 U_g22827 ( .A(I29610), .ZN(g22827) );
INV_X32 U_I29613 ( .A(g21053), .ZN(I29613) );
INV_X32 U_g22828 ( .A(I29613), .ZN(g22828) );
INV_X32 U_g22829 ( .A(g21214), .ZN(g22829) );
INV_X32 U_I29619 ( .A(g21054), .ZN(I29619) );
INV_X32 U_g22832 ( .A(I29619), .ZN(g22832) );
INV_X32 U_I29622 ( .A(g21055), .ZN(I29622) );
INV_X32 U_g22833 ( .A(I29622), .ZN(g22833) );
INV_X32 U_I29625 ( .A(g21056), .ZN(I29625) );
INV_X32 U_g22834 ( .A(I29625), .ZN(g22834) );
INV_X32 U_I29629 ( .A(g21060), .ZN(I29629) );
INV_X32 U_g22836 ( .A(I29629), .ZN(g22836) );
INV_X32 U_I29632 ( .A(g21061), .ZN(I29632) );
INV_X32 U_g22837 ( .A(I29632), .ZN(g22837) );
INV_X32 U_I29635 ( .A(g21062), .ZN(I29635) );
INV_X32 U_g22838 ( .A(I29635), .ZN(g22838) );
INV_X32 U_I29638 ( .A(g21063), .ZN(I29638) );
INV_X32 U_g22839 ( .A(I29638), .ZN(g22839) );
INV_X32 U_I29641 ( .A(g20825), .ZN(I29641) );
INV_X32 U_g22840 ( .A(I29641), .ZN(g22840) );
INV_X32 U_g22843 ( .A(g21889), .ZN(g22843) );
INV_X32 U_g22847 ( .A(g21643), .ZN(g22847) );
INV_X32 U_I29653 ( .A(g21746), .ZN(I29653) );
INV_X32 U_g22852 ( .A(I29653), .ZN(g22852) );
INV_X32 U_I29656 ( .A(g21070), .ZN(I29656) );
INV_X32 U_g22864 ( .A(I29656), .ZN(g22864) );
INV_X32 U_I29660 ( .A(g21071), .ZN(I29660) );
INV_X32 U_g22866 ( .A(I29660), .ZN(g22866) );
INV_X32 U_I29663 ( .A(g21072), .ZN(I29663) );
INV_X32 U_g22867 ( .A(I29663), .ZN(g22867) );
INV_X32 U_g22868 ( .A(g21222), .ZN(g22868) );
INV_X32 U_I29669 ( .A(g21073), .ZN(I29669) );
INV_X32 U_g22871 ( .A(I29669), .ZN(g22871) );
INV_X32 U_I29672 ( .A(g21074), .ZN(I29672) );
INV_X32 U_g22872 ( .A(I29672), .ZN(g22872) );
INV_X32 U_I29675 ( .A(g21075), .ZN(I29675) );
INV_X32 U_g22873 ( .A(I29675), .ZN(g22873) );
INV_X32 U_g22875 ( .A(g21884), .ZN(g22875) );
INV_X32 U_g22882 ( .A(g21674), .ZN(g22882) );
INV_X32 U_I29687 ( .A(g21770), .ZN(I29687) );
INV_X32 U_g22887 ( .A(I29687), .ZN(g22887) );
INV_X32 U_I29690 ( .A(g21080), .ZN(I29690) );
INV_X32 U_g22899 ( .A(I29690), .ZN(g22899) );
INV_X32 U_I29694 ( .A(g21081), .ZN(I29694) );
INV_X32 U_g22901 ( .A(I29694), .ZN(g22901) );
INV_X32 U_I29697 ( .A(g21082), .ZN(I29697) );
INV_X32 U_g22902 ( .A(I29697), .ZN(g22902) );
INV_X32 U_I29700 ( .A(g20700), .ZN(I29700) );
INV_X32 U_g22903 ( .A(I29700), .ZN(g22903) );
INV_X32 U_g22907 ( .A(g21711), .ZN(g22907) );
INV_X32 U_g22917 ( .A(g21703), .ZN(g22917) );
INV_X32 U_I29712 ( .A(g21786), .ZN(I29712) );
INV_X32 U_g22922 ( .A(I29712), .ZN(g22922) );
INV_X32 U_I29715 ( .A(g21094), .ZN(I29715) );
INV_X32 U_g22934 ( .A(I29715), .ZN(g22934) );
INV_X32 U_I29724 ( .A(g21851), .ZN(I29724) );
INV_X32 U_g22945 ( .A(I29724), .ZN(g22945) );
INV_X32 U_I29727 ( .A(g20877), .ZN(I29727) );
INV_X32 U_g22948 ( .A(I29727), .ZN(g22948) );
INV_X32 U_g22949 ( .A(g21665), .ZN(g22949) );
INV_X32 U_g22954 ( .A(g21739), .ZN(g22954) );
INV_X32 U_g22958 ( .A(g21694), .ZN(g22958) );
INV_X32 U_g22962 ( .A(g21763), .ZN(g22962) );
INV_X32 U_g22966 ( .A(g21730), .ZN(g22966) );
INV_X32 U_I29736 ( .A(g20884), .ZN(I29736) );
INV_X32 U_g22970 ( .A(I29736), .ZN(g22970) );
INV_X32 U_g22971 ( .A(g21779), .ZN(g22971) );
INV_X32 U_g22975 ( .A(g21756), .ZN(g22975) );
INV_X32 U_I29741 ( .A(g21346), .ZN(I29741) );
INV_X32 U_g22979 ( .A(I29741), .ZN(g22979) );
INV_X32 U_g22980 ( .A(g21794), .ZN(g22980) );
INV_X32 U_g22986 ( .A(g21382), .ZN(g22986) );
INV_X32 U_g22988 ( .A(g21404), .ZN(g22988) );
INV_X32 U_g22989 ( .A(g21415), .ZN(g22989) );
INV_X32 U_g22991 ( .A(g21429), .ZN(g22991) );
INV_X32 U_g22995 ( .A(g21441), .ZN(g22995) );
INV_X32 U_g22996 ( .A(g21449), .ZN(g22996) );
INV_X32 U_g22998 ( .A(g21458), .ZN(g22998) );
INV_X32 U_g23001 ( .A(g21473), .ZN(g23001) );
INV_X32 U_g23002 ( .A(g21477), .ZN(g23002) );
INV_X32 U_g23006 ( .A(g21483), .ZN(g23006) );
INV_X32 U_g23007 ( .A(g21491), .ZN(g23007) );
INV_X32 U_g23008 ( .A(g21498), .ZN(g23008) );
INV_X32 U_g23012 ( .A(g21505), .ZN(g23012) );
INV_X32 U_g23015 ( .A(g21514), .ZN(g23015) );
INV_X32 U_g23016 ( .A(g21518), .ZN(g23016) );
INV_X32 U_g23020 ( .A(g21524), .ZN(g23020) );
INV_X32 U_g23021 ( .A(g21530), .ZN(g23021) );
INV_X32 U_g23024 ( .A(g21537), .ZN(g23024) );
INV_X32 U_g23028 ( .A(g21541), .ZN(g23028) );
INV_X32 U_g23031 ( .A(g21550), .ZN(g23031) );
INV_X32 U_g23032 ( .A(g21554), .ZN(g23032) );
INV_X32 U_g23036 ( .A(g21558), .ZN(g23036) );
INV_X32 U_g23037 ( .A(g21561), .ZN(g23037) );
INV_X32 U_g23038 ( .A(g21566), .ZN(g23038) );
INV_X32 U_g23041 ( .A(g21573), .ZN(g23041) );
INV_X32 U_g23045 ( .A(g21577), .ZN(g23045) );
INV_X32 U_g23048 ( .A(g21586), .ZN(g23048) );
INV_X32 U_g23049 ( .A(g21590), .ZN(g23049) );
INV_X32 U_I29797 ( .A(g21432), .ZN(I29797) );
INV_X32 U_g23050 ( .A(I29797), .ZN(g23050) );
INV_X32 U_I29802 ( .A(g21435), .ZN(I29802) );
INV_X32 U_g23055 ( .A(I29802), .ZN(g23055) );
INV_X32 U_g23056 ( .A(g21594), .ZN(g23056) );
INV_X32 U_g23057 ( .A(g21599), .ZN(g23057) );
INV_X32 U_g23060 ( .A(g21606), .ZN(g23060) );
INV_X32 U_g23064 ( .A(g21612), .ZN(g23064) );
INV_X32 U_I29812 ( .A(g21467), .ZN(I29812) );
INV_X32 U_g23065 ( .A(I29812), .ZN(g23065) );
INV_X32 U_I29817 ( .A(g21470), .ZN(I29817) );
INV_X32 U_g23068 ( .A(I29817), .ZN(g23068) );
INV_X32 U_g23069 ( .A(g21619), .ZN(g23069) );
INV_X32 U_g23074 ( .A(g21623), .ZN(g23074) );
INV_X32 U_g23075 ( .A(g21628), .ZN(g23075) );
INV_X32 U_I29827 ( .A(g21502), .ZN(I29827) );
INV_X32 U_g23078 ( .A(I29827), .ZN(g23078) );
INV_X32 U_g23079 ( .A(g21640), .ZN(g23079) );
INV_X32 U_g23082 ( .A(g21647), .ZN(g23082) );
INV_X32 U_g23087 ( .A(g21651), .ZN(g23087) );
INV_X32 U_g23088 ( .A(g21655), .ZN(g23088) );
INV_X32 U_I29841 ( .A(g21316), .ZN(I29841) );
INV_X32 U_g23094 ( .A(I29841), .ZN(g23094) );
INV_X32 U_g23095 ( .A(g21671), .ZN(g23095) );
INV_X32 U_g23098 ( .A(g21678), .ZN(g23098) );
INV_X32 U_g23103 ( .A(g21682), .ZN(g23103) );
INV_X32 U_I29852 ( .A(g21331), .ZN(I29852) );
INV_X32 U_g23105 ( .A(I29852), .ZN(g23105) );
INV_X32 U_g23112 ( .A(g21700), .ZN(g23112) );
INV_X32 U_g23115 ( .A(g21708), .ZN(g23115) );
INV_X32 U_I29863 ( .A(g21346), .ZN(I29863) );
INV_X32 U_g23116 ( .A(I29863), .ZN(g23116) );
INV_X32 U_I29872 ( .A(g21364), .ZN(I29872) );
INV_X32 U_g23125 ( .A(I29872), .ZN(g23125) );
INV_X32 U_I29881 ( .A(g21385), .ZN(I29881) );
INV_X32 U_g23134 ( .A(I29881), .ZN(g23134) );
INV_X32 U_g23140 ( .A(g21825), .ZN(g23140) );
INV_X32 U_g23141 ( .A(g21825), .ZN(g23141) );
INV_X32 U_g23142 ( .A(g21825), .ZN(g23142) );
INV_X32 U_g23143 ( .A(g21825), .ZN(g23143) );
INV_X32 U_g23144 ( .A(g21825), .ZN(g23144) );
INV_X32 U_g23145 ( .A(g21825), .ZN(g23145) );
INV_X32 U_g23146 ( .A(g21825), .ZN(g23146) );
INV_X32 U_g23147 ( .A(g21825), .ZN(g23147) );
INV_X32 U_I29897 ( .A(g23116), .ZN(I29897) );
INV_X32 U_g23148 ( .A(I29897), .ZN(g23148) );
INV_X32 U_I29900 ( .A(g23125), .ZN(I29900) );
INV_X32 U_g23149 ( .A(I29900), .ZN(g23149) );
INV_X32 U_I29903 ( .A(g23134), .ZN(I29903) );
INV_X32 U_g23150 ( .A(I29903), .ZN(g23150) );
INV_X32 U_I29906 ( .A(g21967), .ZN(I29906) );
INV_X32 U_g23151 ( .A(I29906), .ZN(g23151) );
INV_X32 U_I29909 ( .A(g23050), .ZN(I29909) );
INV_X32 U_g23152 ( .A(I29909), .ZN(g23152) );
INV_X32 U_I29912 ( .A(g23065), .ZN(I29912) );
INV_X32 U_g23153 ( .A(I29912), .ZN(g23153) );
INV_X32 U_I29915 ( .A(g23055), .ZN(I29915) );
INV_X32 U_g23154 ( .A(I29915), .ZN(g23154) );
INV_X32 U_I29918 ( .A(g23068), .ZN(I29918) );
INV_X32 U_g23155 ( .A(I29918), .ZN(g23155) );
INV_X32 U_I29921 ( .A(g23078), .ZN(I29921) );
INV_X32 U_g23156 ( .A(I29921), .ZN(g23156) );
INV_X32 U_I29924 ( .A(g23094), .ZN(I29924) );
INV_X32 U_g23157 ( .A(I29924), .ZN(g23157) );
INV_X32 U_I29927 ( .A(g23105), .ZN(I29927) );
INV_X32 U_g23158 ( .A(I29927), .ZN(g23158) );
INV_X32 U_I29930 ( .A(g22176), .ZN(I29930) );
INV_X32 U_g23159 ( .A(I29930), .ZN(g23159) );
INV_X32 U_I29933 ( .A(g22082), .ZN(I29933) );
INV_X32 U_g23160 ( .A(I29933), .ZN(g23160) );
INV_X32 U_I29936 ( .A(g22582), .ZN(I29936) );
INV_X32 U_g23161 ( .A(I29936), .ZN(g23161) );
INV_X32 U_I29939 ( .A(g22518), .ZN(I29939) );
INV_X32 U_g23162 ( .A(I29939), .ZN(g23162) );
INV_X32 U_I29942 ( .A(g22548), .ZN(I29942) );
INV_X32 U_g23163 ( .A(I29942), .ZN(g23163) );
INV_X32 U_I29945 ( .A(g22583), .ZN(I29945) );
INV_X32 U_g23164 ( .A(I29945), .ZN(g23164) );
INV_X32 U_I29948 ( .A(g22549), .ZN(I29948) );
INV_X32 U_g23165 ( .A(I29948), .ZN(g23165) );
INV_X32 U_I29951 ( .A(g22584), .ZN(I29951) );
INV_X32 U_g23166 ( .A(I29951), .ZN(g23166) );
INV_X32 U_I29954 ( .A(g22611), .ZN(I29954) );
INV_X32 U_g23167 ( .A(I29954), .ZN(g23167) );
INV_X32 U_I29957 ( .A(g22585), .ZN(I29957) );
INV_X32 U_g23168 ( .A(I29957), .ZN(g23168) );
INV_X32 U_I29960 ( .A(g22612), .ZN(I29960) );
INV_X32 U_g23169 ( .A(I29960), .ZN(g23169) );
INV_X32 U_I29963 ( .A(g22639), .ZN(I29963) );
INV_X32 U_g23170 ( .A(I29963), .ZN(g23170) );
INV_X32 U_I29966 ( .A(g22613), .ZN(I29966) );
INV_X32 U_g23171 ( .A(I29966), .ZN(g23171) );
INV_X32 U_I29969 ( .A(g22640), .ZN(I29969) );
INV_X32 U_g23172 ( .A(I29969), .ZN(g23172) );
INV_X32 U_I29972 ( .A(g22669), .ZN(I29972) );
INV_X32 U_g23173 ( .A(I29972), .ZN(g23173) );
INV_X32 U_I29975 ( .A(g22641), .ZN(I29975) );
INV_X32 U_g23174 ( .A(I29975), .ZN(g23174) );
INV_X32 U_I29978 ( .A(g22670), .ZN(I29978) );
INV_X32 U_g23175 ( .A(I29978), .ZN(g23175) );
INV_X32 U_I29981 ( .A(g22702), .ZN(I29981) );
INV_X32 U_g23176 ( .A(I29981), .ZN(g23176) );
INV_X32 U_I29984 ( .A(g22671), .ZN(I29984) );
INV_X32 U_g23177 ( .A(I29984), .ZN(g23177) );
INV_X32 U_I29987 ( .A(g22703), .ZN(I29987) );
INV_X32 U_g23178 ( .A(I29987), .ZN(g23178) );
INV_X32 U_I29990 ( .A(g22728), .ZN(I29990) );
INV_X32 U_g23179 ( .A(I29990), .ZN(g23179) );
INV_X32 U_I29993 ( .A(g22704), .ZN(I29993) );
INV_X32 U_g23180 ( .A(I29993), .ZN(g23180) );
INV_X32 U_I29996 ( .A(g22729), .ZN(I29996) );
INV_X32 U_g23181 ( .A(I29996), .ZN(g23181) );
INV_X32 U_I29999 ( .A(g22756), .ZN(I29999) );
INV_X32 U_g23182 ( .A(I29999), .ZN(g23182) );
INV_X32 U_I30002 ( .A(g22730), .ZN(I30002) );
INV_X32 U_g23183 ( .A(I30002), .ZN(g23183) );
INV_X32 U_I30005 ( .A(g22757), .ZN(I30005) );
INV_X32 U_g23184 ( .A(I30005), .ZN(g23184) );
INV_X32 U_I30008 ( .A(g22785), .ZN(I30008) );
INV_X32 U_g23185 ( .A(I30008), .ZN(g23185) );
INV_X32 U_I30011 ( .A(g22758), .ZN(I30011) );
INV_X32 U_g23186 ( .A(I30011), .ZN(g23186) );
INV_X32 U_I30014 ( .A(g22786), .ZN(I30014) );
INV_X32 U_g23187 ( .A(I30014), .ZN(g23187) );
INV_X32 U_I30017 ( .A(g22824), .ZN(I30017) );
INV_X32 U_g23188 ( .A(I30017), .ZN(g23188) );
INV_X32 U_I30020 ( .A(g22519), .ZN(I30020) );
INV_X32 U_g23189 ( .A(I30020), .ZN(g23189) );
INV_X32 U_I30023 ( .A(g22550), .ZN(I30023) );
INV_X32 U_g23190 ( .A(I30023), .ZN(g23190) );
INV_X32 U_I30026 ( .A(g22586), .ZN(I30026) );
INV_X32 U_g23191 ( .A(I30026), .ZN(g23191) );
INV_X32 U_I30029 ( .A(g22642), .ZN(I30029) );
INV_X32 U_g23192 ( .A(I30029), .ZN(g23192) );
INV_X32 U_I30032 ( .A(g22672), .ZN(I30032) );
INV_X32 U_g23193 ( .A(I30032), .ZN(g23193) );
INV_X32 U_I30035 ( .A(g22705), .ZN(I30035) );
INV_X32 U_g23194 ( .A(I30035), .ZN(g23194) );
INV_X32 U_I30038 ( .A(g22673), .ZN(I30038) );
INV_X32 U_g23195 ( .A(I30038), .ZN(g23195) );
INV_X32 U_I30041 ( .A(g22706), .ZN(I30041) );
INV_X32 U_g23196 ( .A(I30041), .ZN(g23196) );
INV_X32 U_I30044 ( .A(g22731), .ZN(I30044) );
INV_X32 U_g23197 ( .A(I30044), .ZN(g23197) );
INV_X32 U_I30047 ( .A(g22107), .ZN(I30047) );
INV_X32 U_g23198 ( .A(I30047), .ZN(g23198) );
INV_X32 U_I30050 ( .A(g22619), .ZN(I30050) );
INV_X32 U_g23199 ( .A(I30050), .ZN(g23199) );
INV_X32 U_I30053 ( .A(g22558), .ZN(I30053) );
INV_X32 U_g23200 ( .A(I30053), .ZN(g23200) );
INV_X32 U_I30056 ( .A(g22589), .ZN(I30056) );
INV_X32 U_g23201 ( .A(I30056), .ZN(g23201) );
INV_X32 U_I30059 ( .A(g22620), .ZN(I30059) );
INV_X32 U_g23202 ( .A(I30059), .ZN(g23202) );
INV_X32 U_I30062 ( .A(g22590), .ZN(I30062) );
INV_X32 U_g23203 ( .A(I30062), .ZN(g23203) );
INV_X32 U_I30065 ( .A(g22621), .ZN(I30065) );
INV_X32 U_g23204 ( .A(I30065), .ZN(g23204) );
INV_X32 U_I30068 ( .A(g22647), .ZN(I30068) );
INV_X32 U_g23205 ( .A(I30068), .ZN(g23205) );
INV_X32 U_I30071 ( .A(g22622), .ZN(I30071) );
INV_X32 U_g23206 ( .A(I30071), .ZN(g23206) );
INV_X32 U_I30074 ( .A(g22648), .ZN(I30074) );
INV_X32 U_g23207 ( .A(I30074), .ZN(g23207) );
INV_X32 U_I30077 ( .A(g22675), .ZN(I30077) );
INV_X32 U_g23208 ( .A(I30077), .ZN(g23208) );
INV_X32 U_I30080 ( .A(g22649), .ZN(I30080) );
INV_X32 U_g23209 ( .A(I30080), .ZN(g23209) );
INV_X32 U_I30083 ( .A(g22676), .ZN(I30083) );
INV_X32 U_g23210 ( .A(I30083), .ZN(g23210) );
INV_X32 U_I30086 ( .A(g22709), .ZN(I30086) );
INV_X32 U_g23211 ( .A(I30086), .ZN(g23211) );
INV_X32 U_I30089 ( .A(g22677), .ZN(I30089) );
INV_X32 U_g23212 ( .A(I30089), .ZN(g23212) );
INV_X32 U_I30092 ( .A(g22710), .ZN(I30092) );
INV_X32 U_g23213 ( .A(I30092), .ZN(g23213) );
INV_X32 U_I30095 ( .A(g22733), .ZN(I30095) );
INV_X32 U_g23214 ( .A(I30095), .ZN(g23214) );
INV_X32 U_I30098 ( .A(g22711), .ZN(I30098) );
INV_X32 U_g23215 ( .A(I30098), .ZN(g23215) );
INV_X32 U_I30101 ( .A(g22734), .ZN(I30101) );
INV_X32 U_g23216 ( .A(I30101), .ZN(g23216) );
INV_X32 U_I30104 ( .A(g22760), .ZN(I30104) );
INV_X32 U_g23217 ( .A(I30104), .ZN(g23217) );
INV_X32 U_I30107 ( .A(g22735), .ZN(I30107) );
INV_X32 U_g23218 ( .A(I30107), .ZN(g23218) );
INV_X32 U_I30110 ( .A(g22761), .ZN(I30110) );
INV_X32 U_g23219 ( .A(I30110), .ZN(g23219) );
INV_X32 U_I30113 ( .A(g22790), .ZN(I30113) );
INV_X32 U_g23220 ( .A(I30113), .ZN(g23220) );
INV_X32 U_I30116 ( .A(g22762), .ZN(I30116) );
INV_X32 U_g23221 ( .A(I30116), .ZN(g23221) );
INV_X32 U_I30119 ( .A(g22791), .ZN(I30119) );
INV_X32 U_g23222 ( .A(I30119), .ZN(g23222) );
INV_X32 U_I30122 ( .A(g22827), .ZN(I30122) );
INV_X32 U_g23223 ( .A(I30122), .ZN(g23223) );
INV_X32 U_I30125 ( .A(g22792), .ZN(I30125) );
INV_X32 U_g23224 ( .A(I30125), .ZN(g23224) );
INV_X32 U_I30128 ( .A(g22828), .ZN(I30128) );
INV_X32 U_g23225 ( .A(I30128), .ZN(g23225) );
INV_X32 U_I30131 ( .A(g22864), .ZN(I30131) );
INV_X32 U_g23226 ( .A(I30131), .ZN(g23226) );
INV_X32 U_I30134 ( .A(g22559), .ZN(I30134) );
INV_X32 U_g23227 ( .A(I30134), .ZN(g23227) );
INV_X32 U_I30137 ( .A(g22591), .ZN(I30137) );
INV_X32 U_g23228 ( .A(I30137), .ZN(g23228) );
INV_X32 U_I30140 ( .A(g22623), .ZN(I30140) );
INV_X32 U_g23229 ( .A(I30140), .ZN(g23229) );
INV_X32 U_I30143 ( .A(g22678), .ZN(I30143) );
INV_X32 U_g23230 ( .A(I30143), .ZN(g23230) );
INV_X32 U_I30146 ( .A(g22712), .ZN(I30146) );
INV_X32 U_g23231 ( .A(I30146), .ZN(g23231) );
INV_X32 U_I30149 ( .A(g22736), .ZN(I30149) );
INV_X32 U_g23232 ( .A(I30149), .ZN(g23232) );
INV_X32 U_I30152 ( .A(g22713), .ZN(I30152) );
INV_X32 U_g23233 ( .A(I30152), .ZN(g23233) );
INV_X32 U_I30155 ( .A(g22737), .ZN(I30155) );
INV_X32 U_g23234 ( .A(I30155), .ZN(g23234) );
INV_X32 U_I30158 ( .A(g22763), .ZN(I30158) );
INV_X32 U_g23235 ( .A(I30158), .ZN(g23235) );
INV_X32 U_I30161 ( .A(g22133), .ZN(I30161) );
INV_X32 U_g23236 ( .A(I30161), .ZN(g23236) );
INV_X32 U_I30164 ( .A(g22655), .ZN(I30164) );
INV_X32 U_g23237 ( .A(I30164), .ZN(g23237) );
INV_X32 U_I30167 ( .A(g22598), .ZN(I30167) );
INV_X32 U_g23238 ( .A(I30167), .ZN(g23238) );
INV_X32 U_I30170 ( .A(g22626), .ZN(I30170) );
INV_X32 U_g23239 ( .A(I30170), .ZN(g23239) );
INV_X32 U_I30173 ( .A(g22656), .ZN(I30173) );
INV_X32 U_g23240 ( .A(I30173), .ZN(g23240) );
INV_X32 U_I30176 ( .A(g22627), .ZN(I30176) );
INV_X32 U_g23241 ( .A(I30176), .ZN(g23241) );
INV_X32 U_I30179 ( .A(g22657), .ZN(I30179) );
INV_X32 U_g23242 ( .A(I30179), .ZN(g23242) );
INV_X32 U_I30182 ( .A(g22683), .ZN(I30182) );
INV_X32 U_g23243 ( .A(I30182), .ZN(g23243) );
INV_X32 U_I30185 ( .A(g22658), .ZN(I30185) );
INV_X32 U_g23244 ( .A(I30185), .ZN(g23244) );
INV_X32 U_I30188 ( .A(g22684), .ZN(I30188) );
INV_X32 U_g23245 ( .A(I30188), .ZN(g23245) );
INV_X32 U_I30191 ( .A(g22715), .ZN(I30191) );
INV_X32 U_g23246 ( .A(I30191), .ZN(g23246) );
INV_X32 U_I30194 ( .A(g22685), .ZN(I30194) );
INV_X32 U_g23247 ( .A(I30194), .ZN(g23247) );
INV_X32 U_I30197 ( .A(g22716), .ZN(I30197) );
INV_X32 U_g23248 ( .A(I30197), .ZN(g23248) );
INV_X32 U_I30200 ( .A(g22740), .ZN(I30200) );
INV_X32 U_g23249 ( .A(I30200), .ZN(g23249) );
INV_X32 U_I30203 ( .A(g22717), .ZN(I30203) );
INV_X32 U_g23250 ( .A(I30203), .ZN(g23250) );
INV_X32 U_I30206 ( .A(g22741), .ZN(I30206) );
INV_X32 U_g23251 ( .A(I30206), .ZN(g23251) );
INV_X32 U_I30209 ( .A(g22765), .ZN(I30209) );
INV_X32 U_g23252 ( .A(I30209), .ZN(g23252) );
INV_X32 U_I30212 ( .A(g22742), .ZN(I30212) );
INV_X32 U_g23253 ( .A(I30212), .ZN(g23253) );
INV_X32 U_I30215 ( .A(g22766), .ZN(I30215) );
INV_X32 U_g23254 ( .A(I30215), .ZN(g23254) );
INV_X32 U_I30218 ( .A(g22794), .ZN(I30218) );
INV_X32 U_g23255 ( .A(I30218), .ZN(g23255) );
INV_X32 U_I30221 ( .A(g22767), .ZN(I30221) );
INV_X32 U_g23256 ( .A(I30221), .ZN(g23256) );
INV_X32 U_I30224 ( .A(g22795), .ZN(I30224) );
INV_X32 U_g23257 ( .A(I30224), .ZN(g23257) );
INV_X32 U_I30227 ( .A(g22832), .ZN(I30227) );
INV_X32 U_g23258 ( .A(I30227), .ZN(g23258) );
INV_X32 U_I30230 ( .A(g22796), .ZN(I30230) );
INV_X32 U_g23259 ( .A(I30230), .ZN(g23259) );
INV_X32 U_I30233 ( .A(g22833), .ZN(I30233) );
INV_X32 U_g23260 ( .A(I30233), .ZN(g23260) );
INV_X32 U_I30236 ( .A(g22866), .ZN(I30236) );
INV_X32 U_g23261 ( .A(I30236), .ZN(g23261) );
INV_X32 U_I30239 ( .A(g22834), .ZN(I30239) );
INV_X32 U_g23262 ( .A(I30239), .ZN(g23262) );
INV_X32 U_I30242 ( .A(g22867), .ZN(I30242) );
INV_X32 U_g23263 ( .A(I30242), .ZN(g23263) );
INV_X32 U_I30245 ( .A(g22899), .ZN(I30245) );
INV_X32 U_g23264 ( .A(I30245), .ZN(g23264) );
INV_X32 U_I30248 ( .A(g22599), .ZN(I30248) );
INV_X32 U_g23265 ( .A(I30248), .ZN(g23265) );
INV_X32 U_I30251 ( .A(g22628), .ZN(I30251) );
INV_X32 U_g23266 ( .A(I30251), .ZN(g23266) );
INV_X32 U_I30254 ( .A(g22659), .ZN(I30254) );
INV_X32 U_g23267 ( .A(I30254), .ZN(g23267) );
INV_X32 U_I30257 ( .A(g22718), .ZN(I30257) );
INV_X32 U_g23268 ( .A(I30257), .ZN(g23268) );
INV_X32 U_I30260 ( .A(g22743), .ZN(I30260) );
INV_X32 U_g23269 ( .A(I30260), .ZN(g23269) );
INV_X32 U_I30263 ( .A(g22768), .ZN(I30263) );
INV_X32 U_g23270 ( .A(I30263), .ZN(g23270) );
INV_X32 U_I30266 ( .A(g22744), .ZN(I30266) );
INV_X32 U_g23271 ( .A(I30266), .ZN(g23271) );
INV_X32 U_I30269 ( .A(g22769), .ZN(I30269) );
INV_X32 U_g23272 ( .A(I30269), .ZN(g23272) );
INV_X32 U_I30272 ( .A(g22797), .ZN(I30272) );
INV_X32 U_g23273 ( .A(I30272), .ZN(g23273) );
INV_X32 U_I30275 ( .A(g22156), .ZN(I30275) );
INV_X32 U_g23274 ( .A(I30275), .ZN(g23274) );
INV_X32 U_I30278 ( .A(g22691), .ZN(I30278) );
INV_X32 U_g23275 ( .A(I30278), .ZN(g23275) );
INV_X32 U_I30281 ( .A(g22635), .ZN(I30281) );
INV_X32 U_g23276 ( .A(I30281), .ZN(g23276) );
INV_X32 U_I30284 ( .A(g22662), .ZN(I30284) );
INV_X32 U_g23277 ( .A(I30284), .ZN(g23277) );
INV_X32 U_I30287 ( .A(g22692), .ZN(I30287) );
INV_X32 U_g23278 ( .A(I30287), .ZN(g23278) );
INV_X32 U_I30290 ( .A(g22663), .ZN(I30290) );
INV_X32 U_g23279 ( .A(I30290), .ZN(g23279) );
INV_X32 U_I30293 ( .A(g22693), .ZN(I30293) );
INV_X32 U_g23280 ( .A(I30293), .ZN(g23280) );
INV_X32 U_I30296 ( .A(g22723), .ZN(I30296) );
INV_X32 U_g23281 ( .A(I30296), .ZN(g23281) );
INV_X32 U_I30299 ( .A(g22694), .ZN(I30299) );
INV_X32 U_g23282 ( .A(I30299), .ZN(g23282) );
INV_X32 U_I30302 ( .A(g22724), .ZN(I30302) );
INV_X32 U_g23283 ( .A(I30302), .ZN(g23283) );
INV_X32 U_I30305 ( .A(g22746), .ZN(I30305) );
INV_X32 U_g23284 ( .A(I30305), .ZN(g23284) );
INV_X32 U_I30308 ( .A(g22725), .ZN(I30308) );
INV_X32 U_g23285 ( .A(I30308), .ZN(g23285) );
INV_X32 U_I30311 ( .A(g22747), .ZN(I30311) );
INV_X32 U_g23286 ( .A(I30311), .ZN(g23286) );
INV_X32 U_I30314 ( .A(g22772), .ZN(I30314) );
INV_X32 U_g23287 ( .A(I30314), .ZN(g23287) );
INV_X32 U_I30317 ( .A(g22748), .ZN(I30317) );
INV_X32 U_g23288 ( .A(I30317), .ZN(g23288) );
INV_X32 U_I30320 ( .A(g22773), .ZN(I30320) );
INV_X32 U_g23289 ( .A(I30320), .ZN(g23289) );
INV_X32 U_I30323 ( .A(g22799), .ZN(I30323) );
INV_X32 U_g23290 ( .A(I30323), .ZN(g23290) );
INV_X32 U_I30326 ( .A(g22774), .ZN(I30326) );
INV_X32 U_g23291 ( .A(I30326), .ZN(g23291) );
INV_X32 U_I30329 ( .A(g22800), .ZN(I30329) );
INV_X32 U_g23292 ( .A(I30329), .ZN(g23292) );
INV_X32 U_I30332 ( .A(g22836), .ZN(I30332) );
INV_X32 U_g23293 ( .A(I30332), .ZN(g23293) );
INV_X32 U_I30335 ( .A(g22801), .ZN(I30335) );
INV_X32 U_g23294 ( .A(I30335), .ZN(g23294) );
INV_X32 U_I30338 ( .A(g22837), .ZN(I30338) );
INV_X32 U_g23295 ( .A(I30338), .ZN(g23295) );
INV_X32 U_I30341 ( .A(g22871), .ZN(I30341) );
INV_X32 U_g23296 ( .A(I30341), .ZN(g23296) );
INV_X32 U_I30344 ( .A(g22838), .ZN(I30344) );
INV_X32 U_g23297 ( .A(I30344), .ZN(g23297) );
INV_X32 U_I30347 ( .A(g22872), .ZN(I30347) );
INV_X32 U_g23298 ( .A(I30347), .ZN(g23298) );
INV_X32 U_I30350 ( .A(g22901), .ZN(I30350) );
INV_X32 U_g23299 ( .A(I30350), .ZN(g23299) );
INV_X32 U_I30353 ( .A(g22873), .ZN(I30353) );
INV_X32 U_g23300 ( .A(I30353), .ZN(g23300) );
INV_X32 U_I30356 ( .A(g22902), .ZN(I30356) );
INV_X32 U_g23301 ( .A(I30356), .ZN(g23301) );
INV_X32 U_I30359 ( .A(g22934), .ZN(I30359) );
INV_X32 U_g23302 ( .A(I30359), .ZN(g23302) );
INV_X32 U_I30362 ( .A(g22636), .ZN(I30362) );
INV_X32 U_g23303 ( .A(I30362), .ZN(g23303) );
INV_X32 U_I30365 ( .A(g22664), .ZN(I30365) );
INV_X32 U_g23304 ( .A(I30365), .ZN(g23304) );
INV_X32 U_I30368 ( .A(g22695), .ZN(I30368) );
INV_X32 U_g23305 ( .A(I30368), .ZN(g23305) );
INV_X32 U_I30371 ( .A(g22749), .ZN(I30371) );
INV_X32 U_g23306 ( .A(I30371), .ZN(g23306) );
INV_X32 U_I30374 ( .A(g22775), .ZN(I30374) );
INV_X32 U_g23307 ( .A(I30374), .ZN(g23307) );
INV_X32 U_I30377 ( .A(g22802), .ZN(I30377) );
INV_X32 U_g23308 ( .A(I30377), .ZN(g23308) );
INV_X32 U_I30380 ( .A(g22776), .ZN(I30380) );
INV_X32 U_g23309 ( .A(I30380), .ZN(g23309) );
INV_X32 U_I30383 ( .A(g22803), .ZN(I30383) );
INV_X32 U_g23310 ( .A(I30383), .ZN(g23310) );
INV_X32 U_I30386 ( .A(g22839), .ZN(I30386) );
INV_X32 U_g23311 ( .A(I30386), .ZN(g23311) );
INV_X32 U_I30389 ( .A(g22225), .ZN(I30389) );
INV_X32 U_g23312 ( .A(I30389), .ZN(g23312) );
INV_X32 U_I30392 ( .A(g22226), .ZN(I30392) );
INV_X32 U_g23313 ( .A(I30392), .ZN(g23313) );
INV_X32 U_I30395 ( .A(g22253), .ZN(I30395) );
INV_X32 U_g23314 ( .A(I30395), .ZN(g23314) );
INV_X32 U_I30398 ( .A(g22840), .ZN(I30398) );
INV_X32 U_g23315 ( .A(I30398), .ZN(g23315) );
INV_X32 U_I30401 ( .A(g22444), .ZN(I30401) );
INV_X32 U_g23316 ( .A(I30401), .ZN(g23316) );
INV_X32 U_I30404 ( .A(g22948), .ZN(I30404) );
INV_X32 U_g23317 ( .A(I30404), .ZN(g23317) );
INV_X32 U_I30407 ( .A(g22970), .ZN(I30407) );
INV_X32 U_g23318 ( .A(I30407), .ZN(g23318) );
INV_X32 U_g23403 ( .A(g23052), .ZN(g23403) );
INV_X32 U_g23410 ( .A(g23071), .ZN(g23410) );
INV_X32 U_g23415 ( .A(g23084), .ZN(g23415) );
INV_X32 U_g23420 ( .A(g23089), .ZN(g23420) );
INV_X32 U_g23424 ( .A(g23100), .ZN(g23424) );
INV_X32 U_g23429 ( .A(g23107), .ZN(g23429) );
INV_X32 U_g23435 ( .A(g23120), .ZN(g23435) );
INV_X32 U_I30467 ( .A(g23000), .ZN(I30467) );
INV_X32 U_g23438 ( .A(I30467), .ZN(g23438) );
INV_X32 U_I30470 ( .A(g23117), .ZN(I30470) );
INV_X32 U_g23439 ( .A(I30470), .ZN(g23439) );
INV_X32 U_g23441 ( .A(g23129), .ZN(g23441) );
INV_X32 U_g23444 ( .A(g22945), .ZN(g23444) );
INV_X32 U_I30476 ( .A(g22876), .ZN(I30476) );
INV_X32 U_g23448 ( .A(I30476), .ZN(g23448) );
INV_X32 U_I30480 ( .A(g23014), .ZN(I30480) );
INV_X32 U_g23452 ( .A(I30480), .ZN(g23452) );
INV_X32 U_I30483 ( .A(g23126), .ZN(I30483) );
INV_X32 U_g23453 ( .A(I30483), .ZN(g23453) );
INV_X32 U_I30486 ( .A(g23022), .ZN(I30486) );
INV_X32 U_g23454 ( .A(I30486), .ZN(g23454) );
INV_X32 U_I30489 ( .A(g22911), .ZN(I30489) );
INV_X32 U_g23455 ( .A(I30489), .ZN(g23455) );
INV_X32 U_I30493 ( .A(g23030), .ZN(I30493) );
INV_X32 U_g23459 ( .A(I30493), .ZN(g23459) );
INV_X32 U_I30496 ( .A(g23137), .ZN(I30496) );
INV_X32 U_g23460 ( .A(I30496), .ZN(g23460) );
INV_X32 U_I30501 ( .A(g23039), .ZN(I30501) );
INV_X32 U_g23463 ( .A(I30501), .ZN(g23463) );
INV_X32 U_I30504 ( .A(g22936), .ZN(I30504) );
INV_X32 U_g23464 ( .A(I30504), .ZN(g23464) );
INV_X32 U_I30508 ( .A(g23047), .ZN(I30508) );
INV_X32 U_g23468 ( .A(I30508), .ZN(g23468) );
INV_X32 U_I30511 ( .A(g21970), .ZN(I30511) );
INV_X32 U_g23469 ( .A(I30511), .ZN(g23469) );
INV_X32 U_g23470 ( .A(g22188), .ZN(g23470) );
INV_X32 U_I30516 ( .A(g23058), .ZN(I30516) );
INV_X32 U_g23472 ( .A(I30516), .ZN(g23472) );
INV_X32 U_I30519 ( .A(g22942), .ZN(I30519) );
INV_X32 U_g23473 ( .A(I30519), .ZN(g23473) );
INV_X32 U_I30525 ( .A(g23067), .ZN(I30525) );
INV_X32 U_g23481 ( .A(I30525), .ZN(g23481) );
INV_X32 U_g23482 ( .A(g22197), .ZN(g23482) );
INV_X32 U_I30531 ( .A(g23076), .ZN(I30531) );
INV_X32 U_g23485 ( .A(I30531), .ZN(g23485) );
INV_X32 U_I30536 ( .A(g23081), .ZN(I30536) );
INV_X32 U_g23492 ( .A(I30536), .ZN(g23492) );
INV_X32 U_g23493 ( .A(g22203), .ZN(g23493) );
INV_X32 U_I30544 ( .A(g23092), .ZN(I30544) );
INV_X32 U_g23500 ( .A(I30544), .ZN(g23500) );
INV_X32 U_I30547 ( .A(g23093), .ZN(I30547) );
INV_X32 U_g23501 ( .A(I30547), .ZN(g23501) );
INV_X32 U_I30552 ( .A(g23097), .ZN(I30552) );
INV_X32 U_g23508 ( .A(I30552), .ZN(g23508) );
INV_X32 U_g23509 ( .A(g22209), .ZN(g23509) );
INV_X32 U_I30560 ( .A(g23110), .ZN(I30560) );
INV_X32 U_g23516 ( .A(I30560), .ZN(g23516) );
INV_X32 U_I30563 ( .A(g23111), .ZN(I30563) );
INV_X32 U_g23517 ( .A(I30563), .ZN(g23517) );
INV_X32 U_I30568 ( .A(g23114), .ZN(I30568) );
INV_X32 U_g23524 ( .A(I30568), .ZN(g23524) );
INV_X32 U_I30575 ( .A(g23123), .ZN(I30575) );
INV_X32 U_g23531 ( .A(I30575), .ZN(g23531) );
INV_X32 U_I30578 ( .A(g23124), .ZN(I30578) );
INV_X32 U_g23532 ( .A(I30578), .ZN(g23532) );
INV_X32 U_I30586 ( .A(g23132), .ZN(I30586) );
INV_X32 U_g23542 ( .A(I30586), .ZN(g23542) );
INV_X32 U_I30589 ( .A(g23133), .ZN(I30589) );
INV_X32 U_g23543 ( .A(I30589), .ZN(g23543) );
INV_X32 U_I30594 ( .A(g22025), .ZN(I30594) );
INV_X32 U_g23546 ( .A(I30594), .ZN(g23546) );
INV_X32 U_I30598 ( .A(g22027), .ZN(I30598) );
INV_X32 U_g23548 ( .A(I30598), .ZN(g23548) );
INV_X32 U_I30601 ( .A(g22028), .ZN(I30601) );
INV_X32 U_g23549 ( .A(I30601), .ZN(g23549) );
INV_X32 U_I30607 ( .A(g22029), .ZN(I30607) );
INV_X32 U_g23553 ( .A(I30607), .ZN(g23553) );
INV_X32 U_I30611 ( .A(g22030), .ZN(I30611) );
INV_X32 U_g23555 ( .A(I30611), .ZN(g23555) );
INV_X32 U_I30614 ( .A(g22031), .ZN(I30614) );
INV_X32 U_g23556 ( .A(I30614), .ZN(g23556) );
INV_X32 U_I30617 ( .A(g22032), .ZN(I30617) );
INV_X32 U_g23557 ( .A(I30617), .ZN(g23557) );
INV_X32 U_I30623 ( .A(g22033), .ZN(I30623) );
INV_X32 U_g23561 ( .A(I30623), .ZN(g23561) );
INV_X32 U_I30626 ( .A(g22034), .ZN(I30626) );
INV_X32 U_g23562 ( .A(I30626), .ZN(g23562) );
INV_X32 U_I30632 ( .A(g22035), .ZN(I30632) );
INV_X32 U_g23566 ( .A(I30632), .ZN(g23566) );
INV_X32 U_I30636 ( .A(g22037), .ZN(I30636) );
INV_X32 U_g23568 ( .A(I30636), .ZN(g23568) );
INV_X32 U_I30639 ( .A(g22038), .ZN(I30639) );
INV_X32 U_g23569 ( .A(I30639), .ZN(g23569) );
INV_X32 U_I30642 ( .A(g22039), .ZN(I30642) );
INV_X32 U_g23570 ( .A(I30642), .ZN(g23570) );
INV_X32 U_I30648 ( .A(g22040), .ZN(I30648) );
INV_X32 U_g23574 ( .A(I30648), .ZN(g23574) );
INV_X32 U_I30651 ( .A(g22041), .ZN(I30651) );
INV_X32 U_g23575 ( .A(I30651), .ZN(g23575) );
INV_X32 U_I30654 ( .A(g22042), .ZN(I30654) );
INV_X32 U_g23576 ( .A(I30654), .ZN(g23576) );
INV_X32 U_I30660 ( .A(g22043), .ZN(I30660) );
INV_X32 U_g23580 ( .A(I30660), .ZN(g23580) );
INV_X32 U_I30663 ( .A(g22044), .ZN(I30663) );
INV_X32 U_g23581 ( .A(I30663), .ZN(g23581) );
INV_X32 U_I30669 ( .A(g22045), .ZN(I30669) );
INV_X32 U_g23585 ( .A(I30669), .ZN(g23585) );
INV_X32 U_I30673 ( .A(g22047), .ZN(I30673) );
INV_X32 U_g23587 ( .A(I30673), .ZN(g23587) );
INV_X32 U_I30676 ( .A(g22048), .ZN(I30676) );
INV_X32 U_g23588 ( .A(I30676), .ZN(g23588) );
INV_X32 U_I30679 ( .A(g22049), .ZN(I30679) );
INV_X32 U_g23589 ( .A(I30679), .ZN(g23589) );
INV_X32 U_I30686 ( .A(g23136), .ZN(I30686) );
INV_X32 U_g23594 ( .A(I30686), .ZN(g23594) );
INV_X32 U_I30689 ( .A(g22054), .ZN(I30689) );
INV_X32 U_g23595 ( .A(I30689), .ZN(g23595) );
INV_X32 U_I30692 ( .A(g22055), .ZN(I30692) );
INV_X32 U_g23596 ( .A(I30692), .ZN(g23596) );
INV_X32 U_I30695 ( .A(g22056), .ZN(I30695) );
INV_X32 U_g23597 ( .A(I30695), .ZN(g23597) );
INV_X32 U_I30701 ( .A(g22057), .ZN(I30701) );
INV_X32 U_g23601 ( .A(I30701), .ZN(g23601) );
INV_X32 U_I30704 ( .A(g22058), .ZN(I30704) );
INV_X32 U_g23602 ( .A(I30704), .ZN(g23602) );
INV_X32 U_I30707 ( .A(g22059), .ZN(I30707) );
INV_X32 U_g23603 ( .A(I30707), .ZN(g23603) );
INV_X32 U_I30713 ( .A(g22060), .ZN(I30713) );
INV_X32 U_g23607 ( .A(I30713), .ZN(g23607) );
INV_X32 U_I30716 ( .A(g22061), .ZN(I30716) );
INV_X32 U_g23608 ( .A(I30716), .ZN(g23608) );
INV_X32 U_I30722 ( .A(g22063), .ZN(I30722) );
INV_X32 U_g23612 ( .A(I30722), .ZN(g23612) );
INV_X32 U_I30725 ( .A(g22064), .ZN(I30725) );
INV_X32 U_g23613 ( .A(I30725), .ZN(g23613) );
INV_X32 U_I30728 ( .A(g22065), .ZN(I30728) );
INV_X32 U_g23614 ( .A(I30728), .ZN(g23614) );
INV_X32 U_I30735 ( .A(g22066), .ZN(I30735) );
INV_X32 U_g23619 ( .A(I30735), .ZN(g23619) );
INV_X32 U_I30738 ( .A(g22067), .ZN(I30738) );
INV_X32 U_g23620 ( .A(I30738), .ZN(g23620) );
INV_X32 U_I30741 ( .A(g22068), .ZN(I30741) );
INV_X32 U_g23621 ( .A(I30741), .ZN(g23621) );
INV_X32 U_I30748 ( .A(g21969), .ZN(I30748) );
INV_X32 U_g23626 ( .A(I30748), .ZN(g23626) );
INV_X32 U_I30751 ( .A(g22073), .ZN(I30751) );
INV_X32 U_g23627 ( .A(I30751), .ZN(g23627) );
INV_X32 U_I30754 ( .A(g22074), .ZN(I30754) );
INV_X32 U_g23628 ( .A(I30754), .ZN(g23628) );
INV_X32 U_I30757 ( .A(g22075), .ZN(I30757) );
INV_X32 U_g23629 ( .A(I30757), .ZN(g23629) );
INV_X32 U_I30763 ( .A(g22076), .ZN(I30763) );
INV_X32 U_g23633 ( .A(I30763), .ZN(g23633) );
INV_X32 U_I30766 ( .A(g22077), .ZN(I30766) );
INV_X32 U_g23634 ( .A(I30766), .ZN(g23634) );
INV_X32 U_I30769 ( .A(g22078), .ZN(I30769) );
INV_X32 U_g23635 ( .A(I30769), .ZN(g23635) );
INV_X32 U_I30776 ( .A(g22079), .ZN(I30776) );
INV_X32 U_g23640 ( .A(I30776), .ZN(g23640) );
INV_X32 U_I30779 ( .A(g22080), .ZN(I30779) );
INV_X32 U_g23641 ( .A(I30779), .ZN(g23641) );
INV_X32 U_I30782 ( .A(g22081), .ZN(I30782) );
INV_X32 U_g23642 ( .A(I30782), .ZN(g23642) );
INV_X32 U_I30786 ( .A(g22454), .ZN(I30786) );
INV_X32 U_g23644 ( .A(I30786), .ZN(g23644) );
INV_X32 U_I30797 ( .A(g22087), .ZN(I30797) );
INV_X32 U_g23661 ( .A(I30797), .ZN(g23661) );
INV_X32 U_I30800 ( .A(g22088), .ZN(I30800) );
INV_X32 U_g23662 ( .A(I30800), .ZN(g23662) );
INV_X32 U_I30803 ( .A(g22089), .ZN(I30803) );
INV_X32 U_g23663 ( .A(I30803), .ZN(g23663) );
INV_X32 U_I30810 ( .A(g22090), .ZN(I30810) );
INV_X32 U_g23668 ( .A(I30810), .ZN(g23668) );
INV_X32 U_I30813 ( .A(g22091), .ZN(I30813) );
INV_X32 U_g23669 ( .A(I30813), .ZN(g23669) );
INV_X32 U_I30816 ( .A(g22092), .ZN(I30816) );
INV_X32 U_g23670 ( .A(I30816), .ZN(g23670) );
INV_X32 U_I30823 ( .A(g21972), .ZN(I30823) );
INV_X32 U_g23675 ( .A(I30823), .ZN(g23675) );
INV_X32 U_I30826 ( .A(g22097), .ZN(I30826) );
INV_X32 U_g23676 ( .A(I30826), .ZN(g23676) );
INV_X32 U_I30829 ( .A(g22098), .ZN(I30829) );
INV_X32 U_g23677 ( .A(I30829), .ZN(g23677) );
INV_X32 U_I30832 ( .A(g22099), .ZN(I30832) );
INV_X32 U_g23678 ( .A(I30832), .ZN(g23678) );
INV_X32 U_I30838 ( .A(g22100), .ZN(I30838) );
INV_X32 U_g23682 ( .A(I30838), .ZN(g23682) );
INV_X32 U_I30841 ( .A(g22101), .ZN(I30841) );
INV_X32 U_g23683 ( .A(I30841), .ZN(g23683) );
INV_X32 U_I30844 ( .A(g22102), .ZN(I30844) );
INV_X32 U_g23684 ( .A(I30844), .ZN(g23684) );
INV_X32 U_I30847 ( .A(g22103), .ZN(I30847) );
INV_X32 U_g23685 ( .A(I30847), .ZN(g23685) );
INV_X32 U_I30854 ( .A(g22104), .ZN(I30854) );
INV_X32 U_g23690 ( .A(I30854), .ZN(g23690) );
INV_X32 U_I30857 ( .A(g22105), .ZN(I30857) );
INV_X32 U_g23691 ( .A(I30857), .ZN(g23691) );
INV_X32 U_I30860 ( .A(g22106), .ZN(I30860) );
INV_X32 U_g23692 ( .A(I30860), .ZN(g23692) );
INV_X32 U_I30864 ( .A(g22493), .ZN(I30864) );
INV_X32 U_g23694 ( .A(I30864), .ZN(g23694) );
INV_X32 U_I30875 ( .A(g22112), .ZN(I30875) );
INV_X32 U_g23711 ( .A(I30875), .ZN(g23711) );
INV_X32 U_I30878 ( .A(g22113), .ZN(I30878) );
INV_X32 U_g23712 ( .A(I30878), .ZN(g23712) );
INV_X32 U_I30881 ( .A(g22114), .ZN(I30881) );
INV_X32 U_g23713 ( .A(I30881), .ZN(g23713) );
INV_X32 U_I30888 ( .A(g22115), .ZN(I30888) );
INV_X32 U_g23718 ( .A(I30888), .ZN(g23718) );
INV_X32 U_I30891 ( .A(g22116), .ZN(I30891) );
INV_X32 U_g23719 ( .A(I30891), .ZN(g23719) );
INV_X32 U_I30894 ( .A(g22117), .ZN(I30894) );
INV_X32 U_g23720 ( .A(I30894), .ZN(g23720) );
INV_X32 U_I30901 ( .A(g21974), .ZN(I30901) );
INV_X32 U_g23725 ( .A(I30901), .ZN(g23725) );
INV_X32 U_I30905 ( .A(g22122), .ZN(I30905) );
INV_X32 U_g23727 ( .A(I30905), .ZN(g23727) );
INV_X32 U_I30908 ( .A(g22123), .ZN(I30908) );
INV_X32 U_g23728 ( .A(I30908), .ZN(g23728) );
INV_X32 U_I30911 ( .A(g22124), .ZN(I30911) );
INV_X32 U_g23729 ( .A(I30911), .ZN(g23729) );
INV_X32 U_I30914 ( .A(g22125), .ZN(I30914) );
INV_X32 U_g23730 ( .A(I30914), .ZN(g23730) );
INV_X32 U_I30917 ( .A(g22806), .ZN(I30917) );
INV_X32 U_g23731 ( .A(I30917), .ZN(g23731) );
INV_X32 U_I30922 ( .A(g22126), .ZN(I30922) );
INV_X32 U_g23736 ( .A(I30922), .ZN(g23736) );
INV_X32 U_I30925 ( .A(g22127), .ZN(I30925) );
INV_X32 U_g23737 ( .A(I30925), .ZN(g23737) );
INV_X32 U_I30928 ( .A(g22128), .ZN(I30928) );
INV_X32 U_g23738 ( .A(I30928), .ZN(g23738) );
INV_X32 U_I30931 ( .A(g22129), .ZN(I30931) );
INV_X32 U_g23739 ( .A(I30931), .ZN(g23739) );
INV_X32 U_I30938 ( .A(g22130), .ZN(I30938) );
INV_X32 U_g23744 ( .A(I30938), .ZN(g23744) );
INV_X32 U_I30941 ( .A(g22131), .ZN(I30941) );
INV_X32 U_g23745 ( .A(I30941), .ZN(g23745) );
INV_X32 U_I30944 ( .A(g22132), .ZN(I30944) );
INV_X32 U_g23746 ( .A(I30944), .ZN(g23746) );
INV_X32 U_I30948 ( .A(g22536), .ZN(I30948) );
INV_X32 U_g23748 ( .A(I30948), .ZN(g23748) );
INV_X32 U_I30959 ( .A(g22138), .ZN(I30959) );
INV_X32 U_g23765 ( .A(I30959), .ZN(g23765) );
INV_X32 U_I30962 ( .A(g22139), .ZN(I30962) );
INV_X32 U_g23766 ( .A(I30962), .ZN(g23766) );
INV_X32 U_I30965 ( .A(g22140), .ZN(I30965) );
INV_X32 U_g23767 ( .A(I30965), .ZN(g23767) );
INV_X32 U_I30973 ( .A(g22141), .ZN(I30973) );
INV_X32 U_g23773 ( .A(I30973), .ZN(g23773) );
INV_X32 U_I30976 ( .A(g22142), .ZN(I30976) );
INV_X32 U_g23774 ( .A(I30976), .ZN(g23774) );
INV_X32 U_I30979 ( .A(g22143), .ZN(I30979) );
INV_X32 U_g23775 ( .A(I30979), .ZN(g23775) );
INV_X32 U_I30985 ( .A(g22992), .ZN(I30985) );
INV_X32 U_g23779 ( .A(I30985), .ZN(g23779) );
INV_X32 U_I30988 ( .A(g22145), .ZN(I30988) );
INV_X32 U_g23782 ( .A(I30988), .ZN(g23782) );
INV_X32 U_I30991 ( .A(g22146), .ZN(I30991) );
INV_X32 U_g23783 ( .A(I30991), .ZN(g23783) );
INV_X32 U_I30994 ( .A(g22147), .ZN(I30994) );
INV_X32 U_g23784 ( .A(I30994), .ZN(g23784) );
INV_X32 U_I30997 ( .A(g22148), .ZN(I30997) );
INV_X32 U_g23785 ( .A(I30997), .ZN(g23785) );
INV_X32 U_I31000 ( .A(g22847), .ZN(I31000) );
INV_X32 U_g23786 ( .A(I31000), .ZN(g23786) );
INV_X32 U_I31005 ( .A(g22149), .ZN(I31005) );
INV_X32 U_g23791 ( .A(I31005), .ZN(g23791) );
INV_X32 U_I31008 ( .A(g22150), .ZN(I31008) );
INV_X32 U_g23792 ( .A(I31008), .ZN(g23792) );
INV_X32 U_I31011 ( .A(g22151), .ZN(I31011) );
INV_X32 U_g23793 ( .A(I31011), .ZN(g23793) );
INV_X32 U_I31014 ( .A(g22152), .ZN(I31014) );
INV_X32 U_g23794 ( .A(I31014), .ZN(g23794) );
INV_X32 U_I31021 ( .A(g22153), .ZN(I31021) );
INV_X32 U_g23799 ( .A(I31021), .ZN(g23799) );
INV_X32 U_I31024 ( .A(g22154), .ZN(I31024) );
INV_X32 U_g23800 ( .A(I31024), .ZN(g23800) );
INV_X32 U_I31027 ( .A(g22155), .ZN(I31027) );
INV_X32 U_g23801 ( .A(I31027), .ZN(g23801) );
INV_X32 U_I31031 ( .A(g22576), .ZN(I31031) );
INV_X32 U_g23803 ( .A(I31031), .ZN(g23803) );
INV_X32 U_I31043 ( .A(g22161), .ZN(I31043) );
INV_X32 U_g23821 ( .A(I31043), .ZN(g23821) );
INV_X32 U_I31050 ( .A(g22162), .ZN(I31050) );
INV_X32 U_g23826 ( .A(I31050), .ZN(g23826) );
INV_X32 U_I31053 ( .A(g22163), .ZN(I31053) );
INV_X32 U_g23827 ( .A(I31053), .ZN(g23827) );
INV_X32 U_I31056 ( .A(g22164), .ZN(I31056) );
INV_X32 U_g23828 ( .A(I31056), .ZN(g23828) );
INV_X32 U_I31062 ( .A(g23003), .ZN(I31062) );
INV_X32 U_g23832 ( .A(I31062), .ZN(g23832) );
INV_X32 U_I31065 ( .A(g22166), .ZN(I31065) );
INV_X32 U_g23835 ( .A(I31065), .ZN(g23835) );
INV_X32 U_I31068 ( .A(g22167), .ZN(I31068) );
INV_X32 U_g23836 ( .A(I31068), .ZN(g23836) );
INV_X32 U_I31071 ( .A(g22168), .ZN(I31071) );
INV_X32 U_g23837 ( .A(I31071), .ZN(g23837) );
INV_X32 U_I31074 ( .A(g22169), .ZN(I31074) );
INV_X32 U_g23838 ( .A(I31074), .ZN(g23838) );
INV_X32 U_I31077 ( .A(g22882), .ZN(I31077) );
INV_X32 U_g23839 ( .A(I31077), .ZN(g23839) );
INV_X32 U_I31082 ( .A(g22170), .ZN(I31082) );
INV_X32 U_g23844 ( .A(I31082), .ZN(g23844) );
INV_X32 U_I31085 ( .A(g22171), .ZN(I31085) );
INV_X32 U_g23845 ( .A(I31085), .ZN(g23845) );
INV_X32 U_I31088 ( .A(g22172), .ZN(I31088) );
INV_X32 U_g23846 ( .A(I31088), .ZN(g23846) );
INV_X32 U_I31091 ( .A(g22173), .ZN(I31091) );
INV_X32 U_g23847 ( .A(I31091), .ZN(g23847) );
INV_X32 U_g23853 ( .A(g22300), .ZN(g23853) );
INV_X32 U_I31102 ( .A(g22177), .ZN(I31102) );
INV_X32 U_g23856 ( .A(I31102), .ZN(g23856) );
INV_X32 U_I31109 ( .A(g22178), .ZN(I31109) );
INV_X32 U_g23861 ( .A(I31109), .ZN(g23861) );
INV_X32 U_I31112 ( .A(g22179), .ZN(I31112) );
INV_X32 U_g23862 ( .A(I31112), .ZN(g23862) );
INV_X32 U_I31115 ( .A(g22180), .ZN(I31115) );
INV_X32 U_g23863 ( .A(I31115), .ZN(g23863) );
INV_X32 U_I31121 ( .A(g23017), .ZN(I31121) );
INV_X32 U_g23867 ( .A(I31121), .ZN(g23867) );
INV_X32 U_I31124 ( .A(g22182), .ZN(I31124) );
INV_X32 U_g23870 ( .A(I31124), .ZN(g23870) );
INV_X32 U_I31127 ( .A(g22183), .ZN(I31127) );
INV_X32 U_g23871 ( .A(I31127), .ZN(g23871) );
INV_X32 U_I31130 ( .A(g22184), .ZN(I31130) );
INV_X32 U_g23872 ( .A(I31130), .ZN(g23872) );
INV_X32 U_I31133 ( .A(g22185), .ZN(I31133) );
INV_X32 U_g23873 ( .A(I31133), .ZN(g23873) );
INV_X32 U_I31136 ( .A(g22917), .ZN(I31136) );
INV_X32 U_g23874 ( .A(I31136), .ZN(g23874) );
INV_X32 U_I31141 ( .A(g22777), .ZN(I31141) );
INV_X32 U_g23879 ( .A(I31141), .ZN(g23879) );
INV_X32 U_I31144 ( .A(g22935), .ZN(I31144) );
INV_X32 U_g23882 ( .A(I31144), .ZN(g23882) );
INV_X32 U_g23885 ( .A(g22062), .ZN(g23885) );
INV_X32 U_g23887 ( .A(g22328), .ZN(g23887) );
INV_X32 U_I31152 ( .A(g22191), .ZN(I31152) );
INV_X32 U_g23890 ( .A(I31152), .ZN(g23890) );
INV_X32 U_I31159 ( .A(g22192), .ZN(I31159) );
INV_X32 U_g23895 ( .A(I31159), .ZN(g23895) );
INV_X32 U_I31162 ( .A(g22193), .ZN(I31162) );
INV_X32 U_g23896 ( .A(I31162), .ZN(g23896) );
INV_X32 U_I31165 ( .A(g22194), .ZN(I31165) );
INV_X32 U_g23897 ( .A(I31165), .ZN(g23897) );
INV_X32 U_I31171 ( .A(g23033), .ZN(I31171) );
INV_X32 U_g23901 ( .A(I31171), .ZN(g23901) );
INV_X32 U_g23905 ( .A(g22046), .ZN(g23905) );
INV_X32 U_g23908 ( .A(g22353), .ZN(g23908) );
INV_X32 U_I31181 ( .A(g22200), .ZN(I31181) );
INV_X32 U_g23911 ( .A(I31181), .ZN(g23911) );
INV_X32 U_I31188 ( .A(g21989), .ZN(I31188) );
INV_X32 U_g23916 ( .A(I31188), .ZN(g23916) );
INV_X32 U_g23918 ( .A(g22036), .ZN(g23918) );
INV_X32 U_I31195 ( .A(g22578), .ZN(I31195) );
INV_X32 U_g23923 ( .A(I31195), .ZN(g23923) );
INV_X32 U_g23940 ( .A(g22376), .ZN(g23940) );
INV_X32 U_I31205 ( .A(g22002), .ZN(I31205) );
INV_X32 U_g23943 ( .A(I31205), .ZN(g23943) );
INV_X32 U_I31213 ( .A(g22615), .ZN(I31213) );
INV_X32 U_g23955 ( .A(I31213), .ZN(g23955) );
INV_X32 U_I31226 ( .A(g22651), .ZN(I31226) );
INV_X32 U_g23984 ( .A(I31226), .ZN(g23984) );
INV_X32 U_I31232 ( .A(g22026), .ZN(I31232) );
INV_X32 U_g24000 ( .A(I31232), .ZN(g24000) );
INV_X32 U_I31235 ( .A(g22218), .ZN(I31235) );
INV_X32 U_g24001 ( .A(I31235), .ZN(g24001) );
INV_X32 U_I31244 ( .A(g22687), .ZN(I31244) );
INV_X32 U_g24014 ( .A(I31244), .ZN(g24014) );
INV_X32 U_I31250 ( .A(g22953), .ZN(I31250) );
INV_X32 U_g24030 ( .A(I31250), .ZN(g24030) );
INV_X32 U_I31253 ( .A(g22231), .ZN(I31253) );
INV_X32 U_g24033 ( .A(I31253), .ZN(g24033) );
INV_X32 U_I31257 ( .A(g22234), .ZN(I31257) );
INV_X32 U_g24035 ( .A(I31257), .ZN(g24035) );
INV_X32 U_g24047 ( .A(g23023), .ZN(g24047) );
INV_X32 U_I31266 ( .A(g22242), .ZN(I31266) );
INV_X32 U_g24051 ( .A(I31266), .ZN(g24051) );
INV_X32 U_I31270 ( .A(g22247), .ZN(I31270) );
INV_X32 U_g24053 ( .A(I31270), .ZN(g24053) );
INV_X32 U_I31274 ( .A(g22249), .ZN(I31274) );
INV_X32 U_g24055 ( .A(I31274), .ZN(g24055) );
INV_X32 U_g24060 ( .A(g23040), .ZN(g24060) );
INV_X32 U_I31282 ( .A(g22263), .ZN(I31282) );
INV_X32 U_g24064 ( .A(I31282), .ZN(g24064) );
INV_X32 U_I31286 ( .A(g22267), .ZN(I31286) );
INV_X32 U_g24066 ( .A(I31286), .ZN(g24066) );
INV_X32 U_I31290 ( .A(g22269), .ZN(I31290) );
INV_X32 U_g24068 ( .A(I31290), .ZN(g24068) );
INV_X32 U_g24073 ( .A(g23059), .ZN(g24073) );
INV_X32 U_I31298 ( .A(g22280), .ZN(I31298) );
INV_X32 U_g24077 ( .A(I31298), .ZN(g24077) );
INV_X32 U_I31302 ( .A(g22284), .ZN(I31302) );
INV_X32 U_g24079 ( .A(I31302), .ZN(g24079) );
INV_X32 U_g24084 ( .A(g23077), .ZN(g24084) );
INV_X32 U_I31310 ( .A(g22299), .ZN(I31310) );
INV_X32 U_g24088 ( .A(I31310), .ZN(g24088) );
INV_X32 U_g24094 ( .A(g22339), .ZN(g24094) );
INV_X32 U_g24095 ( .A(g22362), .ZN(g24095) );
INV_X32 U_g24096 ( .A(g22405), .ZN(g24096) );
INV_X32 U_g24097 ( .A(g22382), .ZN(g24097) );
INV_X32 U_g24098 ( .A(g22409), .ZN(g24098) );
INV_X32 U_g24099 ( .A(g22412), .ZN(g24099) );
INV_X32 U_g24101 ( .A(g22415), .ZN(g24101) );
INV_X32 U_g24102 ( .A(g22418), .ZN(g24102) );
INV_X32 U_g24103 ( .A(g22397), .ZN(g24103) );
INV_X32 U_g24104 ( .A(g22422), .ZN(g24104) );
INV_X32 U_g24105 ( .A(g22425), .ZN(g24105) );
INV_X32 U_g24106 ( .A(g22428), .ZN(g24106) );
INV_X32 U_g24107 ( .A(g22431), .ZN(g24107) );
INV_X32 U_g24108 ( .A(g22434), .ZN(g24108) );
INV_X32 U_g24110 ( .A(g22437), .ZN(g24110) );
INV_X32 U_g24111 ( .A(g22440), .ZN(g24111) );
INV_X32 U_g24112 ( .A(g22445), .ZN(g24112) );
INV_X32 U_g24113 ( .A(g22448), .ZN(g24113) );
INV_X32 U_g24114 ( .A(g22451), .ZN(g24114) );
INV_X32 U_g24115 ( .A(g22381), .ZN(g24115) );
INV_X32 U_g24121 ( .A(g22455), .ZN(g24121) );
INV_X32 U_g24122 ( .A(g22458), .ZN(g24122) );
INV_X32 U_g24123 ( .A(g22461), .ZN(g24123) );
INV_X32 U_g24124 ( .A(g22464), .ZN(g24124) );
INV_X32 U_g24125 ( .A(g22467), .ZN(g24125) );
INV_X32 U_g24127 ( .A(g22470), .ZN(g24127) );
INV_X32 U_g24128 ( .A(g22473), .ZN(g24128) );
INV_X32 U_g24129 ( .A(g22477), .ZN(g24129) );
INV_X32 U_g24130 ( .A(g22480), .ZN(g24130) );
INV_X32 U_g24131 ( .A(g22484), .ZN(g24131) );
INV_X32 U_g24132 ( .A(g22487), .ZN(g24132) );
INV_X32 U_g24133 ( .A(g22490), .ZN(g24133) );
INV_X32 U_g24134 ( .A(g22396), .ZN(g24134) );
INV_X32 U_g24140 ( .A(g22494), .ZN(g24140) );
INV_X32 U_g24141 ( .A(g22497), .ZN(g24141) );
INV_X32 U_g24142 ( .A(g22500), .ZN(g24142) );
INV_X32 U_g24143 ( .A(g22503), .ZN(g24143) );
INV_X32 U_g24144 ( .A(g22506), .ZN(g24144) );
INV_X32 U_g24146 ( .A(g22509), .ZN(g24146) );
INV_X32 U_g24147 ( .A(g22512), .ZN(g24147) );
INV_X32 U_g24148 ( .A(g22520), .ZN(g24148) );
INV_X32 U_g24149 ( .A(g22523), .ZN(g24149) );
INV_X32 U_g24150 ( .A(g22527), .ZN(g24150) );
INV_X32 U_g24151 ( .A(g22530), .ZN(g24151) );
INV_X32 U_g24152 ( .A(g22533), .ZN(g24152) );
INV_X32 U_g24153 ( .A(g22399), .ZN(g24153) );
INV_X32 U_g24159 ( .A(g22537), .ZN(g24159) );
INV_X32 U_g24160 ( .A(g22540), .ZN(g24160) );
INV_X32 U_g24161 ( .A(g22543), .ZN(g24161) );
INV_X32 U_g24162 ( .A(g22552), .ZN(g24162) );
INV_X32 U_g24163 ( .A(g22560), .ZN(g24163) );
INV_X32 U_g24164 ( .A(g22563), .ZN(g24164) );
INV_X32 U_g24165 ( .A(g22567), .ZN(g24165) );
INV_X32 U_g24166 ( .A(g22570), .ZN(g24166) );
INV_X32 U_g24167 ( .A(g22573), .ZN(g24167) );
INV_X32 U_g24168 ( .A(g22400), .ZN(g24168) );
INV_X32 U_g24175 ( .A(g22592), .ZN(g24175) );
INV_X32 U_g24176 ( .A(g22600), .ZN(g24176) );
INV_X32 U_g24177 ( .A(g22603), .ZN(g24177) );
INV_X32 U_g24180 ( .A(g22629), .ZN(g24180) );
INV_X32 U_I31387 ( .A(g22811), .ZN(I31387) );
INV_X32 U_g24183 ( .A(I31387), .ZN(g24183) );
INV_X32 U_g24210 ( .A(g22696), .ZN(g24210) );
INV_X32 U_g24220 ( .A(g22750), .ZN(g24220) );
INV_X32 U_I31417 ( .A(g22578), .ZN(I31417) );
INV_X32 U_g24233 ( .A(I31417), .ZN(g24233) );
INV_X32 U_I31426 ( .A(g22615), .ZN(I31426) );
INV_X32 U_g24240 ( .A(I31426), .ZN(g24240) );
INV_X32 U_I31436 ( .A(g22651), .ZN(I31436) );
INV_X32 U_g24248 ( .A(I31436), .ZN(g24248) );
INV_X32 U_g24251 ( .A(g22903), .ZN(g24251) );
INV_X32 U_I31445 ( .A(g22687), .ZN(I31445) );
INV_X32 U_g24255 ( .A(I31445), .ZN(g24255) );
INV_X32 U_I31451 ( .A(g23682), .ZN(I31451) );
INV_X32 U_g24259 ( .A(I31451), .ZN(g24259) );
INV_X32 U_I31454 ( .A(g23727), .ZN(I31454) );
INV_X32 U_g24260 ( .A(I31454), .ZN(g24260) );
INV_X32 U_I31457 ( .A(g23773), .ZN(I31457) );
INV_X32 U_g24261 ( .A(I31457), .ZN(g24261) );
INV_X32 U_I31460 ( .A(g23728), .ZN(I31460) );
INV_X32 U_g24262 ( .A(I31460), .ZN(g24262) );
INV_X32 U_I31463 ( .A(g23774), .ZN(I31463) );
INV_X32 U_g24263 ( .A(I31463), .ZN(g24263) );
INV_X32 U_I31466 ( .A(g23821), .ZN(I31466) );
INV_X32 U_g24264 ( .A(I31466), .ZN(g24264) );
INV_X32 U_I31469 ( .A(g23546), .ZN(I31469) );
INV_X32 U_g24265 ( .A(I31469), .ZN(g24265) );
INV_X32 U_I31472 ( .A(g23548), .ZN(I31472) );
INV_X32 U_g24266 ( .A(I31472), .ZN(g24266) );
INV_X32 U_I31475 ( .A(g23555), .ZN(I31475) );
INV_X32 U_g24267 ( .A(I31475), .ZN(g24267) );
INV_X32 U_I31478 ( .A(g23549), .ZN(I31478) );
INV_X32 U_g24268 ( .A(I31478), .ZN(g24268) );
INV_X32 U_I31481 ( .A(g23556), .ZN(I31481) );
INV_X32 U_g24269 ( .A(I31481), .ZN(g24269) );
INV_X32 U_I31484 ( .A(g23568), .ZN(I31484) );
INV_X32 U_g24270 ( .A(I31484), .ZN(g24270) );
INV_X32 U_I31487 ( .A(g23557), .ZN(I31487) );
INV_X32 U_g24271 ( .A(I31487), .ZN(g24271) );
INV_X32 U_I31490 ( .A(g23569), .ZN(I31490) );
INV_X32 U_g24272 ( .A(I31490), .ZN(g24272) );
INV_X32 U_I31493 ( .A(g23587), .ZN(I31493) );
INV_X32 U_g24273 ( .A(I31493), .ZN(g24273) );
INV_X32 U_I31496 ( .A(g23570), .ZN(I31496) );
INV_X32 U_g24274 ( .A(I31496), .ZN(g24274) );
INV_X32 U_I31499 ( .A(g23588), .ZN(I31499) );
INV_X32 U_g24275 ( .A(I31499), .ZN(g24275) );
INV_X32 U_I31502 ( .A(g23612), .ZN(I31502) );
INV_X32 U_g24276 ( .A(I31502), .ZN(g24276) );
INV_X32 U_I31505 ( .A(g23589), .ZN(I31505) );
INV_X32 U_g24277 ( .A(I31505), .ZN(g24277) );
INV_X32 U_I31508 ( .A(g23613), .ZN(I31508) );
INV_X32 U_g24278 ( .A(I31508), .ZN(g24278) );
INV_X32 U_I31511 ( .A(g23640), .ZN(I31511) );
INV_X32 U_g24279 ( .A(I31511), .ZN(g24279) );
INV_X32 U_I31514 ( .A(g23614), .ZN(I31514) );
INV_X32 U_g24280 ( .A(I31514), .ZN(g24280) );
INV_X32 U_I31517 ( .A(g23641), .ZN(I31517) );
INV_X32 U_g24281 ( .A(I31517), .ZN(g24281) );
INV_X32 U_I31520 ( .A(g23683), .ZN(I31520) );
INV_X32 U_g24282 ( .A(I31520), .ZN(g24282) );
INV_X32 U_I31523 ( .A(g23642), .ZN(I31523) );
INV_X32 U_g24283 ( .A(I31523), .ZN(g24283) );
INV_X32 U_I31526 ( .A(g23684), .ZN(I31526) );
INV_X32 U_g24284 ( .A(I31526), .ZN(g24284) );
INV_X32 U_I31529 ( .A(g23729), .ZN(I31529) );
INV_X32 U_g24285 ( .A(I31529), .ZN(g24285) );
INV_X32 U_I31532 ( .A(g23685), .ZN(I31532) );
INV_X32 U_g24286 ( .A(I31532), .ZN(g24286) );
INV_X32 U_I31535 ( .A(g23730), .ZN(I31535) );
INV_X32 U_g24287 ( .A(I31535), .ZN(g24287) );
INV_X32 U_I31538 ( .A(g23775), .ZN(I31538) );
INV_X32 U_g24288 ( .A(I31538), .ZN(g24288) );
INV_X32 U_I31541 ( .A(g23500), .ZN(I31541) );
INV_X32 U_g24289 ( .A(I31541), .ZN(g24289) );
INV_X32 U_I31544 ( .A(g23438), .ZN(I31544) );
INV_X32 U_g24290 ( .A(I31544), .ZN(g24290) );
INV_X32 U_I31547 ( .A(g23454), .ZN(I31547) );
INV_X32 U_g24291 ( .A(I31547), .ZN(g24291) );
INV_X32 U_I31550 ( .A(g23481), .ZN(I31550) );
INV_X32 U_g24292 ( .A(I31550), .ZN(g24292) );
INV_X32 U_I31553 ( .A(g23501), .ZN(I31553) );
INV_X32 U_g24293 ( .A(I31553), .ZN(g24293) );
INV_X32 U_I31556 ( .A(g23439), .ZN(I31556) );
INV_X32 U_g24294 ( .A(I31556), .ZN(g24294) );
INV_X32 U_I31559 ( .A(g24233), .ZN(I31559) );
INV_X32 U_g24295 ( .A(I31559), .ZN(g24295) );
INV_X32 U_I31562 ( .A(g23594), .ZN(I31562) );
INV_X32 U_g24296 ( .A(I31562), .ZN(g24296) );
INV_X32 U_I31565 ( .A(g24001), .ZN(I31565) );
INV_X32 U_g24297 ( .A(I31565), .ZN(g24297) );
INV_X32 U_I31568 ( .A(g24033), .ZN(I31568) );
INV_X32 U_g24298 ( .A(I31568), .ZN(g24298) );
INV_X32 U_I31571 ( .A(g24051), .ZN(I31571) );
INV_X32 U_g24299 ( .A(I31571), .ZN(g24299) );
INV_X32 U_I31574 ( .A(g23736), .ZN(I31574) );
INV_X32 U_g24300 ( .A(I31574), .ZN(g24300) );
INV_X32 U_I31577 ( .A(g23782), .ZN(I31577) );
INV_X32 U_g24301 ( .A(I31577), .ZN(g24301) );
INV_X32 U_I31580 ( .A(g23826), .ZN(I31580) );
INV_X32 U_g24302 ( .A(I31580), .ZN(g24302) );
INV_X32 U_I31583 ( .A(g23783), .ZN(I31583) );
INV_X32 U_g24303 ( .A(I31583), .ZN(g24303) );
INV_X32 U_I31586 ( .A(g23827), .ZN(I31586) );
INV_X32 U_g24304 ( .A(I31586), .ZN(g24304) );
INV_X32 U_I31589 ( .A(g23856), .ZN(I31589) );
INV_X32 U_g24305 ( .A(I31589), .ZN(g24305) );
INV_X32 U_I31592 ( .A(g23553), .ZN(I31592) );
INV_X32 U_g24306 ( .A(I31592), .ZN(g24306) );
INV_X32 U_I31595 ( .A(g23561), .ZN(I31595) );
INV_X32 U_g24307 ( .A(I31595), .ZN(g24307) );
INV_X32 U_I31598 ( .A(g23574), .ZN(I31598) );
INV_X32 U_g24308 ( .A(I31598), .ZN(g24308) );
INV_X32 U_I31601 ( .A(g23562), .ZN(I31601) );
INV_X32 U_g24309 ( .A(I31601), .ZN(g24309) );
INV_X32 U_I31604 ( .A(g23575), .ZN(I31604) );
INV_X32 U_g24310 ( .A(I31604), .ZN(g24310) );
INV_X32 U_I31607 ( .A(g23595), .ZN(I31607) );
INV_X32 U_g24311 ( .A(I31607), .ZN(g24311) );
INV_X32 U_I31610 ( .A(g23576), .ZN(I31610) );
INV_X32 U_g24312 ( .A(I31610), .ZN(g24312) );
INV_X32 U_I31613 ( .A(g23596), .ZN(I31613) );
INV_X32 U_g24313 ( .A(I31613), .ZN(g24313) );
INV_X32 U_I31616 ( .A(g23619), .ZN(I31616) );
INV_X32 U_g24314 ( .A(I31616), .ZN(g24314) );
INV_X32 U_I31619 ( .A(g23597), .ZN(I31619) );
INV_X32 U_g24315 ( .A(I31619), .ZN(g24315) );
INV_X32 U_I31622 ( .A(g23620), .ZN(I31622) );
INV_X32 U_g24316 ( .A(I31622), .ZN(g24316) );
INV_X32 U_I31625 ( .A(g23661), .ZN(I31625) );
INV_X32 U_g24317 ( .A(I31625), .ZN(g24317) );
INV_X32 U_I31628 ( .A(g23621), .ZN(I31628) );
INV_X32 U_g24318 ( .A(I31628), .ZN(g24318) );
INV_X32 U_I31631 ( .A(g23662), .ZN(I31631) );
INV_X32 U_g24319 ( .A(I31631), .ZN(g24319) );
INV_X32 U_I31634 ( .A(g23690), .ZN(I31634) );
INV_X32 U_g24320 ( .A(I31634), .ZN(g24320) );
INV_X32 U_I31637 ( .A(g23663), .ZN(I31637) );
INV_X32 U_g24321 ( .A(I31637), .ZN(g24321) );
INV_X32 U_I31640 ( .A(g23691), .ZN(I31640) );
INV_X32 U_g24322 ( .A(I31640), .ZN(g24322) );
INV_X32 U_I31643 ( .A(g23737), .ZN(I31643) );
INV_X32 U_g24323 ( .A(I31643), .ZN(g24323) );
INV_X32 U_I31646 ( .A(g23692), .ZN(I31646) );
INV_X32 U_g24324 ( .A(I31646), .ZN(g24324) );
INV_X32 U_I31649 ( .A(g23738), .ZN(I31649) );
INV_X32 U_g24325 ( .A(I31649), .ZN(g24325) );
INV_X32 U_I31652 ( .A(g23784), .ZN(I31652) );
INV_X32 U_g24326 ( .A(I31652), .ZN(g24326) );
INV_X32 U_I31655 ( .A(g23739), .ZN(I31655) );
INV_X32 U_g24327 ( .A(I31655), .ZN(g24327) );
INV_X32 U_I31658 ( .A(g23785), .ZN(I31658) );
INV_X32 U_g24328 ( .A(I31658), .ZN(g24328) );
INV_X32 U_I31661 ( .A(g23828), .ZN(I31661) );
INV_X32 U_g24329 ( .A(I31661), .ZN(g24329) );
INV_X32 U_I31664 ( .A(g23516), .ZN(I31664) );
INV_X32 U_g24330 ( .A(I31664), .ZN(g24330) );
INV_X32 U_I31667 ( .A(g23452), .ZN(I31667) );
INV_X32 U_g24331 ( .A(I31667), .ZN(g24331) );
INV_X32 U_I31670 ( .A(g23463), .ZN(I31670) );
INV_X32 U_g24332 ( .A(I31670), .ZN(g24332) );
INV_X32 U_I31673 ( .A(g23492), .ZN(I31673) );
INV_X32 U_g24333 ( .A(I31673), .ZN(g24333) );
INV_X32 U_I31676 ( .A(g23517), .ZN(I31676) );
INV_X32 U_g24334 ( .A(I31676), .ZN(g24334) );
INV_X32 U_I31679 ( .A(g23453), .ZN(I31679) );
INV_X32 U_g24335 ( .A(I31679), .ZN(g24335) );
INV_X32 U_I31682 ( .A(g24240), .ZN(I31682) );
INV_X32 U_g24336 ( .A(I31682), .ZN(g24336) );
INV_X32 U_I31685 ( .A(g23626), .ZN(I31685) );
INV_X32 U_g24337 ( .A(I31685), .ZN(g24337) );
INV_X32 U_I31688 ( .A(g24035), .ZN(I31688) );
INV_X32 U_g24338 ( .A(I31688), .ZN(g24338) );
INV_X32 U_I31691 ( .A(g24053), .ZN(I31691) );
INV_X32 U_g24339 ( .A(I31691), .ZN(g24339) );
INV_X32 U_I31694 ( .A(g24064), .ZN(I31694) );
INV_X32 U_g24340 ( .A(I31694), .ZN(g24340) );
INV_X32 U_I31697 ( .A(g23791), .ZN(I31697) );
INV_X32 U_g24341 ( .A(I31697), .ZN(g24341) );
INV_X32 U_I31700 ( .A(g23835), .ZN(I31700) );
INV_X32 U_g24342 ( .A(I31700), .ZN(g24342) );
INV_X32 U_I31703 ( .A(g23861), .ZN(I31703) );
INV_X32 U_g24343 ( .A(I31703), .ZN(g24343) );
INV_X32 U_I31706 ( .A(g23836), .ZN(I31706) );
INV_X32 U_g24344 ( .A(I31706), .ZN(g24344) );
INV_X32 U_I31709 ( .A(g23862), .ZN(I31709) );
INV_X32 U_g24345 ( .A(I31709), .ZN(g24345) );
INV_X32 U_I31712 ( .A(g23890), .ZN(I31712) );
INV_X32 U_g24346 ( .A(I31712), .ZN(g24346) );
INV_X32 U_I31715 ( .A(g23566), .ZN(I31715) );
INV_X32 U_g24347 ( .A(I31715), .ZN(g24347) );
INV_X32 U_I31718 ( .A(g23580), .ZN(I31718) );
INV_X32 U_g24348 ( .A(I31718), .ZN(g24348) );
INV_X32 U_I31721 ( .A(g23601), .ZN(I31721) );
INV_X32 U_g24349 ( .A(I31721), .ZN(g24349) );
INV_X32 U_I31724 ( .A(g23581), .ZN(I31724) );
INV_X32 U_g24350 ( .A(I31724), .ZN(g24350) );
INV_X32 U_I31727 ( .A(g23602), .ZN(I31727) );
INV_X32 U_g24351 ( .A(I31727), .ZN(g24351) );
INV_X32 U_I31730 ( .A(g23627), .ZN(I31730) );
INV_X32 U_g24352 ( .A(I31730), .ZN(g24352) );
INV_X32 U_I31733 ( .A(g23603), .ZN(I31733) );
INV_X32 U_g24353 ( .A(I31733), .ZN(g24353) );
INV_X32 U_I31736 ( .A(g23628), .ZN(I31736) );
INV_X32 U_g24354 ( .A(I31736), .ZN(g24354) );
INV_X32 U_I31739 ( .A(g23668), .ZN(I31739) );
INV_X32 U_g24355 ( .A(I31739), .ZN(g24355) );
INV_X32 U_I31742 ( .A(g23629), .ZN(I31742) );
INV_X32 U_g24356 ( .A(I31742), .ZN(g24356) );
INV_X32 U_I31745 ( .A(g23669), .ZN(I31745) );
INV_X32 U_g24357 ( .A(I31745), .ZN(g24357) );
INV_X32 U_I31748 ( .A(g23711), .ZN(I31748) );
INV_X32 U_g24358 ( .A(I31748), .ZN(g24358) );
INV_X32 U_I31751 ( .A(g23670), .ZN(I31751) );
INV_X32 U_g24359 ( .A(I31751), .ZN(g24359) );
INV_X32 U_I31754 ( .A(g23712), .ZN(I31754) );
INV_X32 U_g24360 ( .A(I31754), .ZN(g24360) );
INV_X32 U_I31757 ( .A(g23744), .ZN(I31757) );
INV_X32 U_g24361 ( .A(I31757), .ZN(g24361) );
INV_X32 U_I31760 ( .A(g23713), .ZN(I31760) );
INV_X32 U_g24362 ( .A(I31760), .ZN(g24362) );
INV_X32 U_I31763 ( .A(g23745), .ZN(I31763) );
INV_X32 U_g24363 ( .A(I31763), .ZN(g24363) );
INV_X32 U_I31766 ( .A(g23792), .ZN(I31766) );
INV_X32 U_g24364 ( .A(I31766), .ZN(g24364) );
INV_X32 U_I31769 ( .A(g23746), .ZN(I31769) );
INV_X32 U_g24365 ( .A(I31769), .ZN(g24365) );
INV_X32 U_I31772 ( .A(g23793), .ZN(I31772) );
INV_X32 U_g24366 ( .A(I31772), .ZN(g24366) );
INV_X32 U_I31775 ( .A(g23837), .ZN(I31775) );
INV_X32 U_g24367 ( .A(I31775), .ZN(g24367) );
INV_X32 U_I31778 ( .A(g23794), .ZN(I31778) );
INV_X32 U_g24368 ( .A(I31778), .ZN(g24368) );
INV_X32 U_I31781 ( .A(g23838), .ZN(I31781) );
INV_X32 U_g24369 ( .A(I31781), .ZN(g24369) );
INV_X32 U_I31784 ( .A(g23863), .ZN(I31784) );
INV_X32 U_g24370 ( .A(I31784), .ZN(g24370) );
INV_X32 U_I31787 ( .A(g23531), .ZN(I31787) );
INV_X32 U_g24371 ( .A(I31787), .ZN(g24371) );
INV_X32 U_I31790 ( .A(g23459), .ZN(I31790) );
INV_X32 U_g24372 ( .A(I31790), .ZN(g24372) );
INV_X32 U_I31793 ( .A(g23472), .ZN(I31793) );
INV_X32 U_g24373 ( .A(I31793), .ZN(g24373) );
INV_X32 U_I31796 ( .A(g23508), .ZN(I31796) );
INV_X32 U_g24374 ( .A(I31796), .ZN(g24374) );
INV_X32 U_I31799 ( .A(g23532), .ZN(I31799) );
INV_X32 U_g24375 ( .A(I31799), .ZN(g24375) );
INV_X32 U_I31802 ( .A(g23460), .ZN(I31802) );
INV_X32 U_g24376 ( .A(I31802), .ZN(g24376) );
INV_X32 U_I31805 ( .A(g24248), .ZN(I31805) );
INV_X32 U_g24377 ( .A(I31805), .ZN(g24377) );
INV_X32 U_I31808 ( .A(g23675), .ZN(I31808) );
INV_X32 U_g24378 ( .A(I31808), .ZN(g24378) );
INV_X32 U_I31811 ( .A(g24055), .ZN(I31811) );
INV_X32 U_g24379 ( .A(I31811), .ZN(g24379) );
INV_X32 U_I31814 ( .A(g24066), .ZN(I31814) );
INV_X32 U_g24380 ( .A(I31814), .ZN(g24380) );
INV_X32 U_I31817 ( .A(g24077), .ZN(I31817) );
INV_X32 U_g24381 ( .A(I31817), .ZN(g24381) );
INV_X32 U_I31820 ( .A(g23844), .ZN(I31820) );
INV_X32 U_g24382 ( .A(I31820), .ZN(g24382) );
INV_X32 U_I31823 ( .A(g23870), .ZN(I31823) );
INV_X32 U_g24383 ( .A(I31823), .ZN(g24383) );
INV_X32 U_I31826 ( .A(g23895), .ZN(I31826) );
INV_X32 U_g24384 ( .A(I31826), .ZN(g24384) );
INV_X32 U_I31829 ( .A(g23871), .ZN(I31829) );
INV_X32 U_g24385 ( .A(I31829), .ZN(g24385) );
INV_X32 U_I31832 ( .A(g23896), .ZN(I31832) );
INV_X32 U_g24386 ( .A(I31832), .ZN(g24386) );
INV_X32 U_I31835 ( .A(g23911), .ZN(I31835) );
INV_X32 U_g24387 ( .A(I31835), .ZN(g24387) );
INV_X32 U_I31838 ( .A(g23585), .ZN(I31838) );
INV_X32 U_g24388 ( .A(I31838), .ZN(g24388) );
INV_X32 U_I31841 ( .A(g23607), .ZN(I31841) );
INV_X32 U_g24389 ( .A(I31841), .ZN(g24389) );
INV_X32 U_I31844 ( .A(g23633), .ZN(I31844) );
INV_X32 U_g24390 ( .A(I31844), .ZN(g24390) );
INV_X32 U_I31847 ( .A(g23608), .ZN(I31847) );
INV_X32 U_g24391 ( .A(I31847), .ZN(g24391) );
INV_X32 U_I31850 ( .A(g23634), .ZN(I31850) );
INV_X32 U_g24392 ( .A(I31850), .ZN(g24392) );
INV_X32 U_I31853 ( .A(g23676), .ZN(I31853) );
INV_X32 U_g24393 ( .A(I31853), .ZN(g24393) );
INV_X32 U_I31856 ( .A(g23635), .ZN(I31856) );
INV_X32 U_g24394 ( .A(I31856), .ZN(g24394) );
INV_X32 U_I31859 ( .A(g23677), .ZN(I31859) );
INV_X32 U_g24395 ( .A(I31859), .ZN(g24395) );
INV_X32 U_I31862 ( .A(g23718), .ZN(I31862) );
INV_X32 U_g24396 ( .A(I31862), .ZN(g24396) );
INV_X32 U_I31865 ( .A(g23678), .ZN(I31865) );
INV_X32 U_g24397 ( .A(I31865), .ZN(g24397) );
INV_X32 U_I31868 ( .A(g23719), .ZN(I31868) );
INV_X32 U_g24398 ( .A(I31868), .ZN(g24398) );
INV_X32 U_I31871 ( .A(g23765), .ZN(I31871) );
INV_X32 U_g24399 ( .A(I31871), .ZN(g24399) );
INV_X32 U_I31874 ( .A(g23720), .ZN(I31874) );
INV_X32 U_g24400 ( .A(I31874), .ZN(g24400) );
INV_X32 U_I31877 ( .A(g23766), .ZN(I31877) );
INV_X32 U_g24401 ( .A(I31877), .ZN(g24401) );
INV_X32 U_I31880 ( .A(g23799), .ZN(I31880) );
INV_X32 U_g24402 ( .A(I31880), .ZN(g24402) );
INV_X32 U_I31883 ( .A(g23767), .ZN(I31883) );
INV_X32 U_g24403 ( .A(I31883), .ZN(g24403) );
INV_X32 U_I31886 ( .A(g23800), .ZN(I31886) );
INV_X32 U_g24404 ( .A(I31886), .ZN(g24404) );
INV_X32 U_I31889 ( .A(g23845), .ZN(I31889) );
INV_X32 U_g24405 ( .A(I31889), .ZN(g24405) );
INV_X32 U_I31892 ( .A(g23801), .ZN(I31892) );
INV_X32 U_g24406 ( .A(I31892), .ZN(g24406) );
INV_X32 U_I31895 ( .A(g23846), .ZN(I31895) );
INV_X32 U_g24407 ( .A(I31895), .ZN(g24407) );
INV_X32 U_I31898 ( .A(g23872), .ZN(I31898) );
INV_X32 U_g24408 ( .A(I31898), .ZN(g24408) );
INV_X32 U_I31901 ( .A(g23847), .ZN(I31901) );
INV_X32 U_g24409 ( .A(I31901), .ZN(g24409) );
INV_X32 U_I31904 ( .A(g23873), .ZN(I31904) );
INV_X32 U_g24410 ( .A(I31904), .ZN(g24410) );
INV_X32 U_I31907 ( .A(g23897), .ZN(I31907) );
INV_X32 U_g24411 ( .A(I31907), .ZN(g24411) );
INV_X32 U_I31910 ( .A(g23542), .ZN(I31910) );
INV_X32 U_g24412 ( .A(I31910), .ZN(g24412) );
INV_X32 U_I31913 ( .A(g23468), .ZN(I31913) );
INV_X32 U_g24413 ( .A(I31913), .ZN(g24413) );
INV_X32 U_I31916 ( .A(g23485), .ZN(I31916) );
INV_X32 U_g24414 ( .A(I31916), .ZN(g24414) );
INV_X32 U_I31919 ( .A(g23524), .ZN(I31919) );
INV_X32 U_g24415 ( .A(I31919), .ZN(g24415) );
INV_X32 U_I31922 ( .A(g23543), .ZN(I31922) );
INV_X32 U_g24416 ( .A(I31922), .ZN(g24416) );
INV_X32 U_I31925 ( .A(g23469), .ZN(I31925) );
INV_X32 U_g24417 ( .A(I31925), .ZN(g24417) );
INV_X32 U_I31928 ( .A(g24255), .ZN(I31928) );
INV_X32 U_g24418 ( .A(I31928), .ZN(g24418) );
INV_X32 U_I31931 ( .A(g23725), .ZN(I31931) );
INV_X32 U_g24419 ( .A(I31931), .ZN(g24419) );
INV_X32 U_I31934 ( .A(g24068), .ZN(I31934) );
INV_X32 U_g24420 ( .A(I31934), .ZN(g24420) );
INV_X32 U_I31937 ( .A(g24079), .ZN(I31937) );
INV_X32 U_g24421 ( .A(I31937), .ZN(g24421) );
INV_X32 U_I31940 ( .A(g24088), .ZN(I31940) );
INV_X32 U_g24422 ( .A(I31940), .ZN(g24422) );
INV_X32 U_I31943 ( .A(g24000), .ZN(I31943) );
INV_X32 U_g24423 ( .A(I31943), .ZN(g24423) );
INV_X32 U_I31946 ( .A(g23916), .ZN(I31946) );
INV_X32 U_g24424 ( .A(I31946), .ZN(g24424) );
INV_X32 U_I31949 ( .A(g23943), .ZN(I31949) );
INV_X32 U_g24425 ( .A(I31949), .ZN(g24425) );
INV_X32 U_g24482 ( .A(g24183), .ZN(g24482) );
INV_X32 U_I32042 ( .A(g23399), .ZN(I32042) );
INV_X32 U_g24518 ( .A(I32042), .ZN(g24518) );
INV_X32 U_I32057 ( .A(g23406), .ZN(I32057) );
INV_X32 U_g24531 ( .A(I32057), .ZN(g24531) );
INV_X32 U_I32067 ( .A(g24174), .ZN(I32067) );
INV_X32 U_g24539 ( .A(I32067), .ZN(g24539) );
INV_X32 U_I32074 ( .A(g23413), .ZN(I32074) );
INV_X32 U_g24544 ( .A(I32074), .ZN(g24544) );
INV_X32 U_I32081 ( .A(g24178), .ZN(I32081) );
INV_X32 U_g24549 ( .A(I32081), .ZN(g24549) );
INV_X32 U_I32085 ( .A(g24179), .ZN(I32085) );
INV_X32 U_g24551 ( .A(I32085), .ZN(g24551) );
INV_X32 U_I32092 ( .A(g23418), .ZN(I32092) );
INV_X32 U_g24556 ( .A(I32092), .ZN(g24556) );
INV_X32 U_I32098 ( .A(g24181), .ZN(I32098) );
INV_X32 U_g24560 ( .A(I32098), .ZN(g24560) );
INV_X32 U_I32102 ( .A(g24182), .ZN(I32102) );
INV_X32 U_g24562 ( .A(I32102), .ZN(g24562) );
INV_X32 U_I32109 ( .A(g24206), .ZN(I32109) );
INV_X32 U_g24567 ( .A(I32109), .ZN(g24567) );
INV_X32 U_I32112 ( .A(g24207), .ZN(I32112) );
INV_X32 U_g24568 ( .A(I32112), .ZN(g24568) );
INV_X32 U_I32116 ( .A(g24208), .ZN(I32116) );
INV_X32 U_g24570 ( .A(I32116), .ZN(g24570) );
INV_X32 U_I32120 ( .A(g24209), .ZN(I32120) );
INV_X32 U_g24572 ( .A(I32120), .ZN(g24572) );
INV_X32 U_I32126 ( .A(g24212), .ZN(I32126) );
INV_X32 U_g24576 ( .A(I32126), .ZN(g24576) );
INV_X32 U_I32129 ( .A(g24213), .ZN(I32129) );
INV_X32 U_g24577 ( .A(I32129), .ZN(g24577) );
INV_X32 U_I32133 ( .A(g24214), .ZN(I32133) );
INV_X32 U_g24579 ( .A(I32133), .ZN(g24579) );
INV_X32 U_I32137 ( .A(g24215), .ZN(I32137) );
INV_X32 U_g24581 ( .A(I32137), .ZN(g24581) );
INV_X32 U_I32140 ( .A(g24216), .ZN(I32140) );
INV_X32 U_g24582 ( .A(I32140), .ZN(g24582) );
INV_X32 U_I32143 ( .A(g24218), .ZN(I32143) );
INV_X32 U_g24583 ( .A(I32143), .ZN(g24583) );
INV_X32 U_I32146 ( .A(g24219), .ZN(I32146) );
INV_X32 U_g24584 ( .A(I32146), .ZN(g24584) );
INV_X32 U_I32150 ( .A(g24222), .ZN(I32150) );
INV_X32 U_g24586 ( .A(I32150), .ZN(g24586) );
INV_X32 U_I32153 ( .A(g24223), .ZN(I32153) );
INV_X32 U_g24587 ( .A(I32153), .ZN(g24587) );
INV_X32 U_I32156 ( .A(g24225), .ZN(I32156) );
INV_X32 U_g24588 ( .A(I32156), .ZN(g24588) );
INV_X32 U_I32159 ( .A(g24226), .ZN(I32159) );
INV_X32 U_g24589 ( .A(I32159), .ZN(g24589) );
INV_X32 U_I32164 ( .A(g24228), .ZN(I32164) );
INV_X32 U_g24592 ( .A(I32164), .ZN(g24592) );
INV_X32 U_I32167 ( .A(g24230), .ZN(I32167) );
INV_X32 U_g24593 ( .A(I32167), .ZN(g24593) );
INV_X32 U_I32170 ( .A(g24231), .ZN(I32170) );
INV_X32 U_g24594 ( .A(I32170), .ZN(g24594) );
INV_X32 U_I32175 ( .A(g24235), .ZN(I32175) );
INV_X32 U_g24597 ( .A(I32175), .ZN(g24597) );
INV_X32 U_I32178 ( .A(g24237), .ZN(I32178) );
INV_X32 U_g24598 ( .A(I32178), .ZN(g24598) );
INV_X32 U_I32181 ( .A(g24238), .ZN(I32181) );
INV_X32 U_g24599 ( .A(I32181), .ZN(g24599) );
INV_X32 U_I32184 ( .A(g23497), .ZN(I32184) );
INV_X32 U_g24600 ( .A(I32184), .ZN(g24600) );
INV_X32 U_I32189 ( .A(g24243), .ZN(I32189) );
INV_X32 U_g24605 ( .A(I32189), .ZN(g24605) );
INV_X32 U_I32193 ( .A(g23513), .ZN(I32193) );
INV_X32 U_g24607 ( .A(I32193), .ZN(g24607) );
INV_X32 U_I32198 ( .A(g24250), .ZN(I32198) );
INV_X32 U_g24612 ( .A(I32198), .ZN(g24612) );
INV_X32 U_I32203 ( .A(g23528), .ZN(I32203) );
INV_X32 U_g24619 ( .A(I32203), .ZN(g24619) );
INV_X32 U_I32210 ( .A(g23539), .ZN(I32210) );
INV_X32 U_g24630 ( .A(I32210), .ZN(g24630) );
INV_X32 U_g24648 ( .A(g23470), .ZN(g24648) );
INV_X32 U_g24668 ( .A(g23482), .ZN(g24668) );
INV_X32 U_g24687 ( .A(g23493), .ZN(g24687) );
INV_X32 U_g24704 ( .A(g23509), .ZN(g24704) );
INV_X32 U_I32248 ( .A(g23919), .ZN(I32248) );
INV_X32 U_g24734 ( .A(I32248), .ZN(g24734) );
INV_X32 U_I32251 ( .A(g23919), .ZN(I32251) );
INV_X32 U_g24735 ( .A(I32251), .ZN(g24735) );
INV_X32 U_I32281 ( .A(g23950), .ZN(I32281) );
INV_X32 U_g24763 ( .A(I32281), .ZN(g24763) );
INV_X32 U_I32320 ( .A(g23979), .ZN(I32320) );
INV_X32 U_g24784 ( .A(I32320), .ZN(g24784) );
INV_X32 U_I32365 ( .A(g24009), .ZN(I32365) );
INV_X32 U_g24805 ( .A(I32365), .ZN(g24805) );
INV_X32 U_g24815 ( .A(g23448), .ZN(g24815) );
INV_X32 U_I32388 ( .A(g23385), .ZN(I32388) );
INV_X32 U_g24816 ( .A(I32388), .ZN(g24816) );
INV_X32 U_I32419 ( .A(g24043), .ZN(I32419) );
INV_X32 U_g24827 ( .A(I32419), .ZN(g24827) );
INV_X32 U_g24834 ( .A(g23455), .ZN(g24834) );
INV_X32 U_I32439 ( .A(g23392), .ZN(I32439) );
INV_X32 U_g24835 ( .A(I32439), .ZN(g24835) );
INV_X32 U_g24850 ( .A(g23464), .ZN(g24850) );
INV_X32 U_I32487 ( .A(g23400), .ZN(I32487) );
INV_X32 U_g24851 ( .A(I32487), .ZN(g24851) );
INV_X32 U_I32506 ( .A(g23324), .ZN(I32506) );
INV_X32 U_g24856 ( .A(I32506), .ZN(g24856) );
INV_X32 U_g24864 ( .A(g23473), .ZN(g24864) );
INV_X32 U_I32535 ( .A(g23407), .ZN(I32535) );
INV_X32 U_g24865 ( .A(I32535), .ZN(g24865) );
INV_X32 U_I32556 ( .A(g23329), .ZN(I32556) );
INV_X32 U_g24872 ( .A(I32556), .ZN(g24872) );
INV_X32 U_I32583 ( .A(g23330), .ZN(I32583) );
INV_X32 U_g24879 ( .A(I32583), .ZN(g24879) );
INV_X32 U_I32604 ( .A(g23339), .ZN(I32604) );
INV_X32 U_g24886 ( .A(I32604), .ZN(g24886) );
INV_X32 U_g24893 ( .A(g23486), .ZN(g24893) );
INV_X32 U_I32642 ( .A(g23348), .ZN(I32642) );
INV_X32 U_g24903 ( .A(I32642), .ZN(g24903) );
INV_X32 U_g24912 ( .A(g23495), .ZN(g24912) );
INV_X32 U_g24916 ( .A(g23502), .ZN(g24916) );
INV_X32 U_g24929 ( .A(g23511), .ZN(g24929) );
INV_X32 U_g24933 ( .A(g23518), .ZN(g24933) );
INV_X32 U_g24939 ( .A(g23660), .ZN(g24939) );
INV_X32 U_g24941 ( .A(g23526), .ZN(g24941) );
INV_X32 U_g24945 ( .A(g23533), .ZN(g24945) );
INV_X32 U_I32704 ( .A(g23357), .ZN(I32704) );
INV_X32 U_g24949 ( .A(I32704), .ZN(g24949) );
INV_X32 U_g24950 ( .A(g23710), .ZN(g24950) );
INV_X32 U_g24952 ( .A(g23537), .ZN(g24952) );
INV_X32 U_I32716 ( .A(g23358), .ZN(I32716) );
INV_X32 U_g24956 ( .A(I32716), .ZN(g24956) );
INV_X32 U_I32719 ( .A(g23359), .ZN(I32719) );
INV_X32 U_g24957 ( .A(I32719), .ZN(g24957) );
INV_X32 U_g24958 ( .A(g23478), .ZN(g24958) );
INV_X32 U_g24962 ( .A(g23764), .ZN(g24962) );
INV_X32 U_g24969 ( .A(g23489), .ZN(g24969) );
INV_X32 U_g24973 ( .A(g23819), .ZN(g24973) );
INV_X32 U_g24982 ( .A(g23505), .ZN(g24982) );
INV_X32 U_g24993 ( .A(g23521), .ZN(g24993) );
INV_X32 U_g25087 ( .A(g23731), .ZN(g25087) );
INV_X32 U_g25094 ( .A(g23779), .ZN(g25094) );
INV_X32 U_g25095 ( .A(g23786), .ZN(g25095) );
INV_X32 U_I32829 ( .A(g24059), .ZN(I32829) );
INV_X32 U_g25103 ( .A(I32829), .ZN(g25103) );
INV_X32 U_g25104 ( .A(g23832), .ZN(g25104) );
INV_X32 U_g25105 ( .A(g23839), .ZN(g25105) );
INV_X32 U_I32835 ( .A(g24072), .ZN(I32835) );
INV_X32 U_g25109 ( .A(I32835), .ZN(g25109) );
INV_X32 U_g25110 ( .A(g23867), .ZN(g25110) );
INV_X32 U_g25111 ( .A(g23874), .ZN(g25111) );
INV_X32 U_g25115 ( .A(g23879), .ZN(g25115) );
INV_X32 U_g25116 ( .A(g23882), .ZN(g25116) );
INV_X32 U_I32844 ( .A(g23644), .ZN(I32844) );
INV_X32 U_g25118 ( .A(I32844), .ZN(g25118) );
INV_X32 U_I32847 ( .A(g24083), .ZN(I32847) );
INV_X32 U_g25119 ( .A(I32847), .ZN(g25119) );
INV_X32 U_g25120 ( .A(g23901), .ZN(g25120) );
INV_X32 U_I32851 ( .A(g23694), .ZN(I32851) );
INV_X32 U_g25121 ( .A(I32851), .ZN(g25121) );
INV_X32 U_I32854 ( .A(g24092), .ZN(I32854) );
INV_X32 U_g25122 ( .A(I32854), .ZN(g25122) );
INV_X32 U_I32857 ( .A(g23748), .ZN(I32857) );
INV_X32 U_g25123 ( .A(I32857), .ZN(g25123) );
INV_X32 U_I32860 ( .A(g23803), .ZN(I32860) );
INV_X32 U_g25124 ( .A(I32860), .ZN(g25124) );
INV_X32 U_g25126 ( .A(g24030), .ZN(g25126) );
INV_X32 U_I32868 ( .A(g25118), .ZN(I32868) );
INV_X32 U_g25130 ( .A(I32868), .ZN(g25130) );
INV_X32 U_I32871 ( .A(g24518), .ZN(I32871) );
INV_X32 U_g25131 ( .A(I32871), .ZN(g25131) );
INV_X32 U_I32874 ( .A(g24539), .ZN(I32874) );
INV_X32 U_g25132 ( .A(I32874), .ZN(g25132) );
INV_X32 U_I32877 ( .A(g24567), .ZN(I32877) );
INV_X32 U_g25133 ( .A(I32877), .ZN(g25133) );
INV_X32 U_I32880 ( .A(g24581), .ZN(I32880) );
INV_X32 U_g25134 ( .A(I32880), .ZN(g25134) );
INV_X32 U_I32883 ( .A(g24592), .ZN(I32883) );
INV_X32 U_g25135 ( .A(I32883), .ZN(g25135) );
INV_X32 U_I32886 ( .A(g24549), .ZN(I32886) );
INV_X32 U_g25136 ( .A(I32886), .ZN(g25136) );
INV_X32 U_I32889 ( .A(g24568), .ZN(I32889) );
INV_X32 U_g25137 ( .A(I32889), .ZN(g25137) );
INV_X32 U_I32892 ( .A(g24582), .ZN(I32892) );
INV_X32 U_g25138 ( .A(I32892), .ZN(g25138) );
INV_X32 U_I32895 ( .A(g24816), .ZN(I32895) );
INV_X32 U_g25139 ( .A(I32895), .ZN(g25139) );
INV_X32 U_I32898 ( .A(g24856), .ZN(I32898) );
INV_X32 U_g25140 ( .A(I32898), .ZN(g25140) );
INV_X32 U_I32901 ( .A(g25121), .ZN(I32901) );
INV_X32 U_g25141 ( .A(I32901), .ZN(g25141) );
INV_X32 U_I32904 ( .A(g24531), .ZN(I32904) );
INV_X32 U_g25142 ( .A(I32904), .ZN(g25142) );
INV_X32 U_I32907 ( .A(g24551), .ZN(I32907) );
INV_X32 U_g25143 ( .A(I32907), .ZN(g25143) );
INV_X32 U_I32910 ( .A(g24576), .ZN(I32910) );
INV_X32 U_g25144 ( .A(I32910), .ZN(g25144) );
INV_X32 U_I32913 ( .A(g24586), .ZN(I32913) );
INV_X32 U_g25145 ( .A(I32913), .ZN(g25145) );
INV_X32 U_I32916 ( .A(g24597), .ZN(I32916) );
INV_X32 U_g25146 ( .A(I32916), .ZN(g25146) );
INV_X32 U_I32919 ( .A(g24560), .ZN(I32919) );
INV_X32 U_g25147 ( .A(I32919), .ZN(g25147) );
INV_X32 U_I32922 ( .A(g24577), .ZN(I32922) );
INV_X32 U_g25148 ( .A(I32922), .ZN(g25148) );
INV_X32 U_I32925 ( .A(g24587), .ZN(I32925) );
INV_X32 U_g25149 ( .A(I32925), .ZN(g25149) );
INV_X32 U_I32928 ( .A(g24835), .ZN(I32928) );
INV_X32 U_g25150 ( .A(I32928), .ZN(g25150) );
INV_X32 U_I32931 ( .A(g24872), .ZN(I32931) );
INV_X32 U_g25151 ( .A(I32931), .ZN(g25151) );
INV_X32 U_I32934 ( .A(g25123), .ZN(I32934) );
INV_X32 U_g25152 ( .A(I32934), .ZN(g25152) );
INV_X32 U_I32937 ( .A(g24544), .ZN(I32937) );
INV_X32 U_g25153 ( .A(I32937), .ZN(g25153) );
INV_X32 U_I32940 ( .A(g24562), .ZN(I32940) );
INV_X32 U_g25154 ( .A(I32940), .ZN(g25154) );
INV_X32 U_I32943 ( .A(g24583), .ZN(I32943) );
INV_X32 U_g25155 ( .A(I32943), .ZN(g25155) );
INV_X32 U_I32946 ( .A(g24593), .ZN(I32946) );
INV_X32 U_g25156 ( .A(I32946), .ZN(g25156) );
INV_X32 U_I32949 ( .A(g24605), .ZN(I32949) );
INV_X32 U_g25157 ( .A(I32949), .ZN(g25157) );
INV_X32 U_I32952 ( .A(g24570), .ZN(I32952) );
INV_X32 U_g25158 ( .A(I32952), .ZN(g25158) );
INV_X32 U_I32955 ( .A(g24584), .ZN(I32955) );
INV_X32 U_g25159 ( .A(I32955), .ZN(g25159) );
INV_X32 U_I32958 ( .A(g24594), .ZN(I32958) );
INV_X32 U_g25160 ( .A(I32958), .ZN(g25160) );
INV_X32 U_I32961 ( .A(g24851), .ZN(I32961) );
INV_X32 U_g25161 ( .A(I32961), .ZN(g25161) );
INV_X32 U_I32964 ( .A(g24886), .ZN(I32964) );
INV_X32 U_g25162 ( .A(I32964), .ZN(g25162) );
INV_X32 U_I32967 ( .A(g25124), .ZN(I32967) );
INV_X32 U_g25163 ( .A(I32967), .ZN(g25163) );
INV_X32 U_I32970 ( .A(g24556), .ZN(I32970) );
INV_X32 U_g25164 ( .A(I32970), .ZN(g25164) );
INV_X32 U_I32973 ( .A(g24572), .ZN(I32973) );
INV_X32 U_g25165 ( .A(I32973), .ZN(g25165) );
INV_X32 U_I32976 ( .A(g24588), .ZN(I32976) );
INV_X32 U_g25166 ( .A(I32976), .ZN(g25166) );
INV_X32 U_I32979 ( .A(g24598), .ZN(I32979) );
INV_X32 U_g25167 ( .A(I32979), .ZN(g25167) );
INV_X32 U_I32982 ( .A(g24612), .ZN(I32982) );
INV_X32 U_g25168 ( .A(I32982), .ZN(g25168) );
INV_X32 U_I32985 ( .A(g24579), .ZN(I32985) );
INV_X32 U_g25169 ( .A(I32985), .ZN(g25169) );
INV_X32 U_I32988 ( .A(g24589), .ZN(I32988) );
INV_X32 U_g25170 ( .A(I32988), .ZN(g25170) );
INV_X32 U_I32991 ( .A(g24599), .ZN(I32991) );
INV_X32 U_g25171 ( .A(I32991), .ZN(g25171) );
INV_X32 U_I32994 ( .A(g24865), .ZN(I32994) );
INV_X32 U_g25172 ( .A(I32994), .ZN(g25172) );
INV_X32 U_I32997 ( .A(g24903), .ZN(I32997) );
INV_X32 U_g25173 ( .A(I32997), .ZN(g25173) );
INV_X32 U_I33000 ( .A(g24949), .ZN(I33000) );
INV_X32 U_g25174 ( .A(I33000), .ZN(g25174) );
INV_X32 U_I33003 ( .A(g24956), .ZN(I33003) );
INV_X32 U_g25175 ( .A(I33003), .ZN(g25175) );
INV_X32 U_I33006 ( .A(g24957), .ZN(I33006) );
INV_X32 U_g25176 ( .A(I33006), .ZN(g25176) );
INV_X32 U_I33009 ( .A(g24879), .ZN(I33009) );
INV_X32 U_g25177 ( .A(I33009), .ZN(g25177) );
INV_X32 U_I33013 ( .A(g25119), .ZN(I33013) );
INV_X32 U_g25179 ( .A(I33013), .ZN(g25179) );
INV_X32 U_I33016 ( .A(g25122), .ZN(I33016) );
INV_X32 U_g25180 ( .A(I33016), .ZN(g25180) );
INV_X32 U_g25274 ( .A(g24912), .ZN(g25274) );
INV_X32 U_g25283 ( .A(g24929), .ZN(g25283) );
INV_X32 U_g25291 ( .A(g24941), .ZN(g25291) );
INV_X32 U_I33128 ( .A(g24975), .ZN(I33128) );
INV_X32 U_g25296 ( .A(I33128), .ZN(g25296) );
INV_X32 U_g25301 ( .A(g24952), .ZN(g25301) );
INV_X32 U_g25305 ( .A(g24880), .ZN(g25305) );
INV_X32 U_I33136 ( .A(g24986), .ZN(I33136) );
INV_X32 U_g25306 ( .A(I33136), .ZN(g25306) );
INV_X32 U_g25313 ( .A(g24868), .ZN(g25313) );
INV_X32 U_g25314 ( .A(g24897), .ZN(g25314) );
INV_X32 U_I33145 ( .A(g24997), .ZN(I33145) );
INV_X32 U_g25315 ( .A(I33145), .ZN(g25315) );
INV_X32 U_g25319 ( .A(g24857), .ZN(g25319) );
INV_X32 U_g25322 ( .A(g24883), .ZN(g25322) );
INV_X32 U_g25323 ( .A(g24920), .ZN(g25323) );
INV_X32 U_I33154 ( .A(g25005), .ZN(I33154) );
INV_X32 U_g25324 ( .A(I33154), .ZN(g25324) );
INV_X32 U_I33157 ( .A(g25027), .ZN(I33157) );
INV_X32 U_g25327 ( .A(I33157), .ZN(g25327) );
INV_X32 U_g25329 ( .A(g24844), .ZN(g25329) );
INV_X32 U_g25330 ( .A(g24873), .ZN(g25330) );
INV_X32 U_g25332 ( .A(g24900), .ZN(g25332) );
INV_X32 U_g25333 ( .A(g24937), .ZN(g25333) );
INV_X32 U_g25335 ( .A(g24832), .ZN(g25335) );
INV_X32 U_I33168 ( .A(g25042), .ZN(I33168) );
INV_X32 U_g25336 ( .A(I33168), .ZN(g25336) );
INV_X32 U_g25338 ( .A(g24860), .ZN(g25338) );
INV_X32 U_g25339 ( .A(g24887), .ZN(g25339) );
INV_X32 U_g25341 ( .A(g24923), .ZN(g25341) );
INV_X32 U_g25347 ( .A(g24817), .ZN(g25347) );
INV_X32 U_g25349 ( .A(g24848), .ZN(g25349) );
INV_X32 U_I33182 ( .A(g25056), .ZN(I33182) );
INV_X32 U_g25350 ( .A(I33182), .ZN(g25350) );
INV_X32 U_g25352 ( .A(g24875), .ZN(g25352) );
INV_X32 U_g25353 ( .A(g24904), .ZN(g25353) );
INV_X32 U_I33188 ( .A(g24814), .ZN(I33188) );
INV_X32 U_g25354 ( .A(I33188), .ZN(g25354) );
INV_X32 U_g25355 ( .A(g24797), .ZN(g25355) );
INV_X32 U_g25361 ( .A(g24837), .ZN(g25361) );
INV_X32 U_g25363 ( .A(g24862), .ZN(g25363) );
INV_X32 U_I33198 ( .A(g25067), .ZN(I33198) );
INV_X32 U_g25364 ( .A(I33198), .ZN(g25364) );
INV_X32 U_g25366 ( .A(g24889), .ZN(g25366) );
INV_X32 U_g25367 ( .A(g24676), .ZN(g25367) );
INV_X32 U_g25368 ( .A(g24778), .ZN(g25368) );
INV_X32 U_I33205 ( .A(g24833), .ZN(I33205) );
INV_X32 U_g25369 ( .A(I33205), .ZN(g25369) );
INV_X32 U_g25370 ( .A(g24820), .ZN(g25370) );
INV_X32 U_g25376 ( .A(g24852), .ZN(g25376) );
INV_X32 U_g25378 ( .A(g24877), .ZN(g25378) );
INV_X32 U_g25379 ( .A(g24893), .ZN(g25379) );
INV_X32 U_g25383 ( .A(g24766), .ZN(g25383) );
INV_X32 U_g25384 ( .A(g24695), .ZN(g25384) );
INV_X32 U_g25385 ( .A(g24801), .ZN(g25385) );
INV_X32 U_I33219 ( .A(g24849), .ZN(I33219) );
INV_X32 U_g25386 ( .A(I33219), .ZN(g25386) );
INV_X32 U_g25387 ( .A(g24839), .ZN(g25387) );
INV_X32 U_g25393 ( .A(g24866), .ZN(g25393) );
INV_X32 U_g25394 ( .A(g24753), .ZN(g25394) );
INV_X32 U_g25395 ( .A(g24916), .ZN(g25395) );
INV_X32 U_g25399 ( .A(g24787), .ZN(g25399) );
INV_X32 U_g25400 ( .A(g24712), .ZN(g25400) );
INV_X32 U_g25401 ( .A(g24823), .ZN(g25401) );
INV_X32 U_I33232 ( .A(g24863), .ZN(I33232) );
INV_X32 U_g25402 ( .A(I33232), .ZN(g25402) );
INV_X32 U_g25403 ( .A(g24854), .ZN(g25403) );
INV_X32 U_g25404 ( .A(g24771), .ZN(g25404) );
INV_X32 U_g25405 ( .A(g24933), .ZN(g25405) );
INV_X32 U_g25409 ( .A(g24808), .ZN(g25409) );
INV_X32 U_g25410 ( .A(g24723), .ZN(g25410) );
INV_X32 U_g25411 ( .A(g24842), .ZN(g25411) );
INV_X32 U_g25412 ( .A(g24791), .ZN(g25412) );
INV_X32 U_g25413 ( .A(g24945), .ZN(g25413) );
INV_X32 U_g25417 ( .A(g24830), .ZN(g25417) );
INV_X32 U_g25419 ( .A(g24812), .ZN(g25419) );
INV_X32 U_I33246 ( .A(g24890), .ZN(I33246) );
INV_X32 U_g25420 ( .A(I33246), .ZN(g25420) );
INV_X32 U_I33249 ( .A(g24890), .ZN(I33249) );
INV_X32 U_g25421 ( .A(I33249), .ZN(g25421) );
INV_X32 U_g25422 ( .A(g24958), .ZN(g25422) );
INV_X32 U_g25430 ( .A(g24616), .ZN(g25430) );
INV_X32 U_g25431 ( .A(g24969), .ZN(g25431) );
INV_X32 U_I33257 ( .A(g24909), .ZN(I33257) );
INV_X32 U_g25435 ( .A(I33257), .ZN(g25435) );
INV_X32 U_I33260 ( .A(g24909), .ZN(I33260) );
INV_X32 U_g25436 ( .A(I33260), .ZN(g25436) );
INV_X32 U_g25437 ( .A(g24627), .ZN(g25437) );
INV_X32 U_g25438 ( .A(g24982), .ZN(g25438) );
INV_X32 U_I33265 ( .A(g24925), .ZN(I33265) );
INV_X32 U_g25442 ( .A(I33265), .ZN(g25442) );
INV_X32 U_I33268 ( .A(g24925), .ZN(I33268) );
INV_X32 U_g25443 ( .A(I33268), .ZN(g25443) );
INV_X32 U_g25444 ( .A(g24641), .ZN(g25444) );
INV_X32 U_g25445 ( .A(g24993), .ZN(g25445) );
INV_X32 U_g25449 ( .A(g24660), .ZN(g25449) );
INV_X32 U_I33278 ( .A(g25088), .ZN(I33278) );
INV_X32 U_g25454 ( .A(I33278), .ZN(g25454) );
INV_X32 U_I33282 ( .A(g25096), .ZN(I33282) );
INV_X32 U_g25458 ( .A(I33282), .ZN(g25458) );
INV_X32 U_I33286 ( .A(g24426), .ZN(I33286) );
INV_X32 U_g25462 ( .A(I33286), .ZN(g25462) );
INV_X32 U_I33289 ( .A(g25106), .ZN(I33289) );
INV_X32 U_g25463 ( .A(I33289), .ZN(g25463) );
INV_X32 U_I33293 ( .A(g25008), .ZN(I33293) );
INV_X32 U_g25467 ( .A(I33293), .ZN(g25467) );
INV_X32 U_I33297 ( .A(g24430), .ZN(I33297) );
INV_X32 U_g25471 ( .A(I33297), .ZN(g25471) );
INV_X32 U_I33300 ( .A(g25112), .ZN(I33300) );
INV_X32 U_g25472 ( .A(I33300), .ZN(g25472) );
INV_X32 U_I33304 ( .A(g25004), .ZN(I33304) );
INV_X32 U_g25476 ( .A(I33304), .ZN(g25476) );
INV_X32 U_I33307 ( .A(g25011), .ZN(I33307) );
INV_X32 U_g25479 ( .A(I33307), .ZN(g25479) );
INV_X32 U_I33312 ( .A(g25014), .ZN(I33312) );
INV_X32 U_g25484 ( .A(I33312), .ZN(g25484) );
INV_X32 U_I33316 ( .A(g24434), .ZN(I33316) );
INV_X32 U_g25488 ( .A(I33316), .ZN(g25488) );
INV_X32 U_I33321 ( .A(g24442), .ZN(I33321) );
INV_X32 U_g25493 ( .A(I33321), .ZN(g25493) );
INV_X32 U_I33324 ( .A(g25009), .ZN(I33324) );
INV_X32 U_g25496 ( .A(I33324), .ZN(g25496) );
INV_X32 U_I33327 ( .A(g25017), .ZN(I33327) );
INV_X32 U_g25499 ( .A(I33327), .ZN(g25499) );
INV_X32 U_I33330 ( .A(g25019), .ZN(I33330) );
INV_X32 U_g25502 ( .A(I33330), .ZN(g25502) );
INV_X32 U_I33335 ( .A(g25010), .ZN(I33335) );
INV_X32 U_g25507 ( .A(I33335), .ZN(g25507) );
INV_X32 U_I33338 ( .A(g25021), .ZN(I33338) );
INV_X32 U_g25510 ( .A(I33338), .ZN(g25510) );
INV_X32 U_I33343 ( .A(g25024), .ZN(I33343) );
INV_X32 U_g25515 ( .A(I33343), .ZN(g25515) );
INV_X32 U_I33347 ( .A(g24438), .ZN(I33347) );
INV_X32 U_g25519 ( .A(I33347), .ZN(g25519) );
INV_X32 U_I33352 ( .A(g24443), .ZN(I33352) );
INV_X32 U_g25524 ( .A(I33352), .ZN(g25524) );
INV_X32 U_I33355 ( .A(g25012), .ZN(I33355) );
INV_X32 U_g25527 ( .A(I33355), .ZN(g25527) );
INV_X32 U_I33358 ( .A(g25028), .ZN(I33358) );
INV_X32 U_g25530 ( .A(I33358), .ZN(g25530) );
INV_X32 U_I33361 ( .A(g25013), .ZN(I33361) );
INV_X32 U_g25533 ( .A(I33361), .ZN(g25533) );
INV_X32 U_I33364 ( .A(g25029), .ZN(I33364) );
INV_X32 U_g25536 ( .A(I33364), .ZN(g25536) );
INV_X32 U_I33368 ( .A(g24444), .ZN(I33368) );
INV_X32 U_g25540 ( .A(I33368), .ZN(g25540) );
INV_X32 U_I33371 ( .A(g25015), .ZN(I33371) );
INV_X32 U_g25543 ( .A(I33371), .ZN(g25543) );
INV_X32 U_I33374 ( .A(g25031), .ZN(I33374) );
INV_X32 U_g25546 ( .A(I33374), .ZN(g25546) );
INV_X32 U_I33377 ( .A(g25033), .ZN(I33377) );
INV_X32 U_g25549 ( .A(I33377), .ZN(g25549) );
INV_X32 U_I33382 ( .A(g25016), .ZN(I33382) );
INV_X32 U_g25554 ( .A(I33382), .ZN(g25554) );
INV_X32 U_I33385 ( .A(g25035), .ZN(I33385) );
INV_X32 U_g25557 ( .A(I33385), .ZN(g25557) );
INV_X32 U_I33390 ( .A(g25038), .ZN(I33390) );
INV_X32 U_g25562 ( .A(I33390), .ZN(g25562) );
INV_X32 U_I33396 ( .A(g24447), .ZN(I33396) );
INV_X32 U_g25573 ( .A(I33396), .ZN(g25573) );
INV_X32 U_I33399 ( .A(g25018), .ZN(I33399) );
INV_X32 U_g25576 ( .A(I33399), .ZN(g25576) );
INV_X32 U_I33402 ( .A(g24448), .ZN(I33402) );
INV_X32 U_g25579 ( .A(I33402), .ZN(g25579) );
INV_X32 U_I33405 ( .A(g25020), .ZN(I33405) );
INV_X32 U_g25582 ( .A(I33405), .ZN(g25582) );
INV_X32 U_I33408 ( .A(g25040), .ZN(I33408) );
INV_X32 U_g25585 ( .A(I33408), .ZN(g25585) );
INV_X32 U_I33411 ( .A(g24491), .ZN(I33411) );
INV_X32 U_g25588 ( .A(I33411), .ZN(g25588) );
INV_X32 U_I33415 ( .A(g24449), .ZN(I33415) );
INV_X32 U_g25590 ( .A(I33415), .ZN(g25590) );
INV_X32 U_I33418 ( .A(g25022), .ZN(I33418) );
INV_X32 U_g25593 ( .A(I33418), .ZN(g25593) );
INV_X32 U_I33421 ( .A(g25043), .ZN(I33421) );
INV_X32 U_g25596 ( .A(I33421), .ZN(g25596) );
INV_X32 U_I33424 ( .A(g25023), .ZN(I33424) );
INV_X32 U_g25599 ( .A(I33424), .ZN(g25599) );
INV_X32 U_I33427 ( .A(g25044), .ZN(I33427) );
INV_X32 U_g25602 ( .A(I33427), .ZN(g25602) );
INV_X32 U_I33431 ( .A(g24450), .ZN(I33431) );
INV_X32 U_g25606 ( .A(I33431), .ZN(g25606) );
INV_X32 U_I33434 ( .A(g25025), .ZN(I33434) );
INV_X32 U_g25609 ( .A(I33434), .ZN(g25609) );
INV_X32 U_I33437 ( .A(g25046), .ZN(I33437) );
INV_X32 U_g25612 ( .A(I33437), .ZN(g25612) );
INV_X32 U_I33440 ( .A(g25048), .ZN(I33440) );
INV_X32 U_g25615 ( .A(I33440), .ZN(g25615) );
INV_X32 U_I33445 ( .A(g25026), .ZN(I33445) );
INV_X32 U_g25620 ( .A(I33445), .ZN(g25620) );
INV_X32 U_I33448 ( .A(g25050), .ZN(I33448) );
INV_X32 U_g25623 ( .A(I33448), .ZN(g25623) );
INV_X32 U_g25630 ( .A(g24478), .ZN(g25630) );
INV_X32 U_I33457 ( .A(g24451), .ZN(I33457) );
INV_X32 U_g25634 ( .A(I33457), .ZN(g25634) );
INV_X32 U_I33460 ( .A(g24452), .ZN(I33460) );
INV_X32 U_g25637 ( .A(I33460), .ZN(g25637) );
INV_X32 U_I33463 ( .A(g25030), .ZN(I33463) );
INV_X32 U_g25640 ( .A(I33463), .ZN(g25640) );
INV_X32 U_I33466 ( .A(g25053), .ZN(I33466) );
INV_X32 U_g25643 ( .A(I33466), .ZN(g25643) );
INV_X32 U_I33469 ( .A(g24498), .ZN(I33469) );
INV_X32 U_g25646 ( .A(I33469), .ZN(g25646) );
INV_X32 U_I33472 ( .A(g24499), .ZN(I33472) );
INV_X32 U_g25647 ( .A(I33472), .ZN(g25647) );
INV_X32 U_I33476 ( .A(g24453), .ZN(I33476) );
INV_X32 U_g25652 ( .A(I33476), .ZN(g25652) );
INV_X32 U_I33479 ( .A(g25032), .ZN(I33479) );
INV_X32 U_g25655 ( .A(I33479), .ZN(g25655) );
INV_X32 U_I33482 ( .A(g24454), .ZN(I33482) );
INV_X32 U_g25658 ( .A(I33482), .ZN(g25658) );
INV_X32 U_I33485 ( .A(g25034), .ZN(I33485) );
INV_X32 U_g25661 ( .A(I33485), .ZN(g25661) );
INV_X32 U_I33488 ( .A(g25054), .ZN(I33488) );
INV_X32 U_g25664 ( .A(I33488), .ZN(g25664) );
INV_X32 U_I33491 ( .A(g24501), .ZN(I33491) );
INV_X32 U_g25667 ( .A(I33491), .ZN(g25667) );
INV_X32 U_I33495 ( .A(g24455), .ZN(I33495) );
INV_X32 U_g25669 ( .A(I33495), .ZN(g25669) );
INV_X32 U_I33498 ( .A(g25036), .ZN(I33498) );
INV_X32 U_g25672 ( .A(I33498), .ZN(g25672) );
INV_X32 U_I33501 ( .A(g25057), .ZN(I33501) );
INV_X32 U_g25675 ( .A(I33501), .ZN(g25675) );
INV_X32 U_I33504 ( .A(g25037), .ZN(I33504) );
INV_X32 U_g25678 ( .A(I33504), .ZN(g25678) );
INV_X32 U_I33507 ( .A(g25058), .ZN(I33507) );
INV_X32 U_g25681 ( .A(I33507), .ZN(g25681) );
INV_X32 U_I33511 ( .A(g24456), .ZN(I33511) );
INV_X32 U_g25685 ( .A(I33511), .ZN(g25685) );
INV_X32 U_I33514 ( .A(g25039), .ZN(I33514) );
INV_X32 U_g25688 ( .A(I33514), .ZN(g25688) );
INV_X32 U_I33517 ( .A(g25060), .ZN(I33517) );
INV_X32 U_g25691 ( .A(I33517), .ZN(g25691) );
INV_X32 U_I33520 ( .A(g25062), .ZN(I33520) );
INV_X32 U_g25694 ( .A(I33520), .ZN(g25694) );
INV_X32 U_g25698 ( .A(g24600), .ZN(g25698) );
INV_X32 U_I33526 ( .A(g24457), .ZN(I33526) );
INV_X32 U_g25700 ( .A(I33526), .ZN(g25700) );
INV_X32 U_I33529 ( .A(g25041), .ZN(I33529) );
INV_X32 U_g25703 ( .A(I33529), .ZN(g25703) );
INV_X32 U_I33532 ( .A(g24507), .ZN(I33532) );
INV_X32 U_g25706 ( .A(I33532), .ZN(g25706) );
INV_X32 U_I33535 ( .A(g24508), .ZN(I33535) );
INV_X32 U_g25707 ( .A(I33535), .ZN(g25707) );
INV_X32 U_I33539 ( .A(g24458), .ZN(I33539) );
INV_X32 U_g25711 ( .A(I33539), .ZN(g25711) );
INV_X32 U_I33542 ( .A(g24459), .ZN(I33542) );
INV_X32 U_g25714 ( .A(I33542), .ZN(g25714) );
INV_X32 U_I33545 ( .A(g25045), .ZN(I33545) );
INV_X32 U_g25717 ( .A(I33545), .ZN(g25717) );
INV_X32 U_I33548 ( .A(g25064), .ZN(I33548) );
INV_X32 U_g25720 ( .A(I33548), .ZN(g25720) );
INV_X32 U_I33551 ( .A(g24510), .ZN(I33551) );
INV_X32 U_g25723 ( .A(I33551), .ZN(g25723) );
INV_X32 U_I33554 ( .A(g24511), .ZN(I33554) );
INV_X32 U_g25724 ( .A(I33554), .ZN(g25724) );
INV_X32 U_I33558 ( .A(g24460), .ZN(I33558) );
INV_X32 U_g25729 ( .A(I33558), .ZN(g25729) );
INV_X32 U_I33561 ( .A(g25047), .ZN(I33561) );
INV_X32 U_g25732 ( .A(I33561), .ZN(g25732) );
INV_X32 U_I33564 ( .A(g24461), .ZN(I33564) );
INV_X32 U_g25735 ( .A(I33564), .ZN(g25735) );
INV_X32 U_I33567 ( .A(g25049), .ZN(I33567) );
INV_X32 U_g25738 ( .A(I33567), .ZN(g25738) );
INV_X32 U_I33570 ( .A(g25065), .ZN(I33570) );
INV_X32 U_g25741 ( .A(I33570), .ZN(g25741) );
INV_X32 U_I33573 ( .A(g24513), .ZN(I33573) );
INV_X32 U_g25744 ( .A(I33573), .ZN(g25744) );
INV_X32 U_I33577 ( .A(g24462), .ZN(I33577) );
INV_X32 U_g25746 ( .A(I33577), .ZN(g25746) );
INV_X32 U_I33580 ( .A(g25051), .ZN(I33580) );
INV_X32 U_g25749 ( .A(I33580), .ZN(g25749) );
INV_X32 U_I33583 ( .A(g25068), .ZN(I33583) );
INV_X32 U_g25752 ( .A(I33583), .ZN(g25752) );
INV_X32 U_I33586 ( .A(g25052), .ZN(I33586) );
INV_X32 U_g25755 ( .A(I33586), .ZN(g25755) );
INV_X32 U_I33589 ( .A(g25069), .ZN(I33589) );
INV_X32 U_g25758 ( .A(I33589), .ZN(g25758) );
INV_X32 U_I33593 ( .A(g24445), .ZN(I33593) );
INV_X32 U_g25762 ( .A(I33593), .ZN(g25762) );
INV_X32 U_I33596 ( .A(g24446), .ZN(I33596) );
INV_X32 U_g25763 ( .A(I33596), .ZN(g25763) );
INV_X32 U_I33600 ( .A(g24463), .ZN(I33600) );
INV_X32 U_g25767 ( .A(I33600), .ZN(g25767) );
INV_X32 U_I33603 ( .A(g24519), .ZN(I33603) );
INV_X32 U_g25770 ( .A(I33603), .ZN(g25770) );
INV_X32 U_g25771 ( .A(g24607), .ZN(g25771) );
INV_X32 U_I33608 ( .A(g24464), .ZN(I33608) );
INV_X32 U_g25773 ( .A(I33608), .ZN(g25773) );
INV_X32 U_I33611 ( .A(g25055), .ZN(I33611) );
INV_X32 U_g25776 ( .A(I33611), .ZN(g25776) );
INV_X32 U_I33614 ( .A(g24521), .ZN(I33614) );
INV_X32 U_g25779 ( .A(I33614), .ZN(g25779) );
INV_X32 U_I33617 ( .A(g24522), .ZN(I33617) );
INV_X32 U_g25780 ( .A(I33617), .ZN(g25780) );
INV_X32 U_I33621 ( .A(g24465), .ZN(I33621) );
INV_X32 U_g25784 ( .A(I33621), .ZN(g25784) );
INV_X32 U_I33624 ( .A(g24466), .ZN(I33624) );
INV_X32 U_g25787 ( .A(I33624), .ZN(g25787) );
INV_X32 U_I33627 ( .A(g25059), .ZN(I33627) );
INV_X32 U_g25790 ( .A(I33627), .ZN(g25790) );
INV_X32 U_I33630 ( .A(g25071), .ZN(I33630) );
INV_X32 U_g25793 ( .A(I33630), .ZN(g25793) );
INV_X32 U_I33633 ( .A(g24524), .ZN(I33633) );
INV_X32 U_g25796 ( .A(I33633), .ZN(g25796) );
INV_X32 U_I33636 ( .A(g24525), .ZN(I33636) );
INV_X32 U_g25797 ( .A(I33636), .ZN(g25797) );
INV_X32 U_I33640 ( .A(g24467), .ZN(I33640) );
INV_X32 U_g25802 ( .A(I33640), .ZN(g25802) );
INV_X32 U_I33643 ( .A(g25061), .ZN(I33643) );
INV_X32 U_g25805 ( .A(I33643), .ZN(g25805) );
INV_X32 U_I33646 ( .A(g24468), .ZN(I33646) );
INV_X32 U_g25808 ( .A(I33646), .ZN(g25808) );
INV_X32 U_I33649 ( .A(g25063), .ZN(I33649) );
INV_X32 U_g25811 ( .A(I33649), .ZN(g25811) );
INV_X32 U_I33652 ( .A(g25072), .ZN(I33652) );
INV_X32 U_g25814 ( .A(I33652), .ZN(g25814) );
INV_X32 U_I33655 ( .A(g24527), .ZN(I33655) );
INV_X32 U_g25817 ( .A(I33655), .ZN(g25817) );
INV_X32 U_I33659 ( .A(g24469), .ZN(I33659) );
INV_X32 U_g25821 ( .A(I33659), .ZN(g25821) );
INV_X32 U_I33662 ( .A(g24532), .ZN(I33662) );
INV_X32 U_g25824 ( .A(I33662), .ZN(g25824) );
INV_X32 U_g25825 ( .A(g24619), .ZN(g25825) );
INV_X32 U_I33667 ( .A(g24470), .ZN(I33667) );
INV_X32 U_g25827 ( .A(I33667), .ZN(g25827) );
INV_X32 U_I33670 ( .A(g25066), .ZN(I33670) );
INV_X32 U_g25830 ( .A(I33670), .ZN(g25830) );
INV_X32 U_I33673 ( .A(g24534), .ZN(I33673) );
INV_X32 U_g25833 ( .A(I33673), .ZN(g25833) );
INV_X32 U_I33676 ( .A(g24535), .ZN(I33676) );
INV_X32 U_g25834 ( .A(I33676), .ZN(g25834) );
INV_X32 U_I33680 ( .A(g24471), .ZN(I33680) );
INV_X32 U_g25838 ( .A(I33680), .ZN(g25838) );
INV_X32 U_I33683 ( .A(g24472), .ZN(I33683) );
INV_X32 U_g25841 ( .A(I33683), .ZN(g25841) );
INV_X32 U_I33686 ( .A(g25070), .ZN(I33686) );
INV_X32 U_g25844 ( .A(I33686), .ZN(g25844) );
INV_X32 U_I33689 ( .A(g25074), .ZN(I33689) );
INV_X32 U_g25847 ( .A(I33689), .ZN(g25847) );
INV_X32 U_I33692 ( .A(g24537), .ZN(I33692) );
INV_X32 U_g25850 ( .A(I33692), .ZN(g25850) );
INV_X32 U_I33695 ( .A(g24538), .ZN(I33695) );
INV_X32 U_g25851 ( .A(I33695), .ZN(g25851) );
INV_X32 U_I33700 ( .A(g24474), .ZN(I33700) );
INV_X32 U_g25856 ( .A(I33700), .ZN(g25856) );
INV_X32 U_I33703 ( .A(g24545), .ZN(I33703) );
INV_X32 U_g25859 ( .A(I33703), .ZN(g25859) );
INV_X32 U_g25860 ( .A(g24630), .ZN(g25860) );
INV_X32 U_I33708 ( .A(g24475), .ZN(I33708) );
INV_X32 U_g25862 ( .A(I33708), .ZN(g25862) );
INV_X32 U_I33711 ( .A(g25073), .ZN(I33711) );
INV_X32 U_g25865 ( .A(I33711), .ZN(g25865) );
INV_X32 U_I33714 ( .A(g24547), .ZN(I33714) );
INV_X32 U_g25868 ( .A(I33714), .ZN(g25868) );
INV_X32 U_I33717 ( .A(g24548), .ZN(I33717) );
INV_X32 U_g25869 ( .A(I33717), .ZN(g25869) );
INV_X32 U_I33723 ( .A(g24477), .ZN(I33723) );
INV_X32 U_g25877 ( .A(I33723), .ZN(g25877) );
INV_X32 U_I33726 ( .A(g24557), .ZN(I33726) );
INV_X32 U_g25880 ( .A(I33726), .ZN(g25880) );
INV_X32 U_I33732 ( .A(g24473), .ZN(I33732) );
INV_X32 U_g25886 ( .A(I33732), .ZN(g25886) );
INV_X32 U_I33737 ( .A(g24476), .ZN(I33737) );
INV_X32 U_g25891 ( .A(I33737), .ZN(g25891) );
INV_X32 U_g25895 ( .A(g24939), .ZN(g25895) );
INV_X32 U_g25899 ( .A(g24928), .ZN(g25899) );
INV_X32 U_g25903 ( .A(g24950), .ZN(g25903) );
INV_X32 U_g25907 ( .A(g24940), .ZN(g25907) );
INV_X32 U_g25911 ( .A(g24962), .ZN(g25911) );
INV_X32 U_g25915 ( .A(g24951), .ZN(g25915) );
INV_X32 U_g25919 ( .A(g24973), .ZN(g25919) );
INV_X32 U_g25923 ( .A(g24963), .ZN(g25923) );
INV_X32 U_g25937 ( .A(g24763), .ZN(g25937) );
INV_X32 U_g25939 ( .A(g24784), .ZN(g25939) );
INV_X32 U_g25942 ( .A(g24805), .ZN(g25942) );
INV_X32 U_g25945 ( .A(g24827), .ZN(g25945) );
INV_X32 U_g25952 ( .A(g24735), .ZN(g25952) );
INV_X32 U_I33790 ( .A(g25103), .ZN(I33790) );
INV_X32 U_g25976 ( .A(I33790), .ZN(g25976) );
INV_X32 U_I33798 ( .A(g25109), .ZN(I33798) );
INV_X32 U_g25982 ( .A(I33798), .ZN(g25982) );
INV_X32 U_I33801 ( .A(g25327), .ZN(I33801) );
INV_X32 U_g25983 ( .A(I33801), .ZN(g25983) );
INV_X32 U_I33804 ( .A(g25976), .ZN(I33804) );
INV_X32 U_g25984 ( .A(I33804), .ZN(g25984) );
INV_X32 U_I33807 ( .A(g25588), .ZN(I33807) );
INV_X32 U_g25985 ( .A(I33807), .ZN(g25985) );
INV_X32 U_I33810 ( .A(g25646), .ZN(I33810) );
INV_X32 U_g25986 ( .A(I33810), .ZN(g25986) );
INV_X32 U_I33813 ( .A(g25706), .ZN(I33813) );
INV_X32 U_g25987 ( .A(I33813), .ZN(g25987) );
INV_X32 U_I33816 ( .A(g25647), .ZN(I33816) );
INV_X32 U_g25988 ( .A(I33816), .ZN(g25988) );
INV_X32 U_I33819 ( .A(g25707), .ZN(I33819) );
INV_X32 U_g25989 ( .A(I33819), .ZN(g25989) );
INV_X32 U_I33822 ( .A(g25770), .ZN(I33822) );
INV_X32 U_g25990 ( .A(I33822), .ZN(g25990) );
INV_X32 U_I33825 ( .A(g25462), .ZN(I33825) );
INV_X32 U_g25991 ( .A(I33825), .ZN(g25991) );
INV_X32 U_I33828 ( .A(g25336), .ZN(I33828) );
INV_X32 U_g25992 ( .A(I33828), .ZN(g25992) );
INV_X32 U_I33831 ( .A(g25982), .ZN(I33831) );
INV_X32 U_g25993 ( .A(I33831), .ZN(g25993) );
INV_X32 U_I33834 ( .A(g25667), .ZN(I33834) );
INV_X32 U_g25994 ( .A(I33834), .ZN(g25994) );
INV_X32 U_I33837 ( .A(g25723), .ZN(I33837) );
INV_X32 U_g25995 ( .A(I33837), .ZN(g25995) );
INV_X32 U_I33840 ( .A(g25779), .ZN(I33840) );
INV_X32 U_g25996 ( .A(I33840), .ZN(g25996) );
INV_X32 U_I33843 ( .A(g25724), .ZN(I33843) );
INV_X32 U_g25997 ( .A(I33843), .ZN(g25997) );
INV_X32 U_I33846 ( .A(g25780), .ZN(I33846) );
INV_X32 U_g25998 ( .A(I33846), .ZN(g25998) );
INV_X32 U_I33849 ( .A(g25824), .ZN(I33849) );
INV_X32 U_g25999 ( .A(I33849), .ZN(g25999) );
INV_X32 U_I33852 ( .A(g25471), .ZN(I33852) );
INV_X32 U_g26000 ( .A(I33852), .ZN(g26000) );
INV_X32 U_I33855 ( .A(g25350), .ZN(I33855) );
INV_X32 U_g26001 ( .A(I33855), .ZN(g26001) );
INV_X32 U_I33858 ( .A(g25179), .ZN(I33858) );
INV_X32 U_g26002 ( .A(I33858), .ZN(g26002) );
INV_X32 U_I33861 ( .A(g25744), .ZN(I33861) );
INV_X32 U_g26003 ( .A(I33861), .ZN(g26003) );
INV_X32 U_I33864 ( .A(g25796), .ZN(I33864) );
INV_X32 U_g26004 ( .A(I33864), .ZN(g26004) );
INV_X32 U_I33867 ( .A(g25833), .ZN(I33867) );
INV_X32 U_g26005 ( .A(I33867), .ZN(g26005) );
INV_X32 U_I33870 ( .A(g25797), .ZN(I33870) );
INV_X32 U_g26006 ( .A(I33870), .ZN(g26006) );
INV_X32 U_I33873 ( .A(g25834), .ZN(I33873) );
INV_X32 U_g26007 ( .A(I33873), .ZN(g26007) );
INV_X32 U_I33876 ( .A(g25859), .ZN(I33876) );
INV_X32 U_g26008 ( .A(I33876), .ZN(g26008) );
INV_X32 U_I33879 ( .A(g25488), .ZN(I33879) );
INV_X32 U_g26009 ( .A(I33879), .ZN(g26009) );
INV_X32 U_I33882 ( .A(g25364), .ZN(I33882) );
INV_X32 U_g26010 ( .A(I33882), .ZN(g26010) );
INV_X32 U_I33885 ( .A(g25180), .ZN(I33885) );
INV_X32 U_g26011 ( .A(I33885), .ZN(g26011) );
INV_X32 U_I33888 ( .A(g25817), .ZN(I33888) );
INV_X32 U_g26012 ( .A(I33888), .ZN(g26012) );
INV_X32 U_I33891 ( .A(g25850), .ZN(I33891) );
INV_X32 U_g26013 ( .A(I33891), .ZN(g26013) );
INV_X32 U_I33894 ( .A(g25868), .ZN(I33894) );
INV_X32 U_g26014 ( .A(I33894), .ZN(g26014) );
INV_X32 U_I33897 ( .A(g25851), .ZN(I33897) );
INV_X32 U_g26015 ( .A(I33897), .ZN(g26015) );
INV_X32 U_I33900 ( .A(g25869), .ZN(I33900) );
INV_X32 U_g26016 ( .A(I33900), .ZN(g26016) );
INV_X32 U_I33903 ( .A(g25880), .ZN(I33903) );
INV_X32 U_g26017 ( .A(I33903), .ZN(g26017) );
INV_X32 U_I33906 ( .A(g25519), .ZN(I33906) );
INV_X32 U_g26018 ( .A(I33906), .ZN(g26018) );
INV_X32 U_I33909 ( .A(g25886), .ZN(I33909) );
INV_X32 U_g26019 ( .A(I33909), .ZN(g26019) );
INV_X32 U_I33912 ( .A(g25891), .ZN(I33912) );
INV_X32 U_g26020 ( .A(I33912), .ZN(g26020) );
INV_X32 U_I33915 ( .A(g25762), .ZN(I33915) );
INV_X32 U_g26021 ( .A(I33915), .ZN(g26021) );
INV_X32 U_I33918 ( .A(g25763), .ZN(I33918) );
INV_X32 U_g26022 ( .A(I33918), .ZN(g26022) );
INV_X32 U_I33954 ( .A(g25343), .ZN(I33954) );
INV_X32 U_g26056 ( .A(I33954), .ZN(g26056) );
INV_X32 U_I33961 ( .A(g25357), .ZN(I33961) );
INV_X32 U_g26063 ( .A(I33961), .ZN(g26063) );
INV_X32 U_I33968 ( .A(g25372), .ZN(I33968) );
INV_X32 U_g26070 ( .A(I33968), .ZN(g26070) );
INV_X32 U_I33974 ( .A(g25389), .ZN(I33974) );
INV_X32 U_g26076 ( .A(I33974), .ZN(g26076) );
INV_X32 U_I33984 ( .A(g25932), .ZN(I33984) );
INV_X32 U_g26086 ( .A(I33984), .ZN(g26086) );
INV_X32 U_I33990 ( .A(g25870), .ZN(I33990) );
INV_X32 U_g26092 ( .A(I33990), .ZN(g26092) );
INV_X32 U_I33995 ( .A(g25935), .ZN(I33995) );
INV_X32 U_g26102 ( .A(I33995), .ZN(g26102) );
INV_X32 U_I33999 ( .A(g25490), .ZN(I33999) );
INV_X32 U_g26104 ( .A(I33999), .ZN(g26104) );
INV_X32 U_I34002 ( .A(g25490), .ZN(I34002) );
INV_X32 U_g26105 ( .A(I34002), .ZN(g26105) );
INV_X32 U_I34009 ( .A(g25882), .ZN(I34009) );
INV_X32 U_g26114 ( .A(I34009), .ZN(g26114) );
INV_X32 U_I34012 ( .A(g25938), .ZN(I34012) );
INV_X32 U_g26118 ( .A(I34012), .ZN(g26118) );
INV_X32 U_I34017 ( .A(g25887), .ZN(I34017) );
INV_X32 U_g26121 ( .A(I34017), .ZN(g26121) );
INV_X32 U_I34020 ( .A(g25940), .ZN(I34020) );
INV_X32 U_g26125 ( .A(I34020), .ZN(g26125) );
INV_X32 U_I34026 ( .A(g25892), .ZN(I34026) );
INV_X32 U_g26131 ( .A(I34026), .ZN(g26131) );
INV_X32 U_I34029 ( .A(g25520), .ZN(I34029) );
INV_X32 U_g26135 ( .A(I34029), .ZN(g26135) );
INV_X32 U_I34032 ( .A(g25520), .ZN(I34032) );
INV_X32 U_g26136 ( .A(I34032), .ZN(g26136) );
INV_X32 U_I34041 ( .A(g25566), .ZN(I34041) );
INV_X32 U_g26149 ( .A(I34041), .ZN(g26149) );
INV_X32 U_I34044 ( .A(g25566), .ZN(I34044) );
INV_X32 U_g26150 ( .A(I34044), .ZN(g26150) );
INV_X32 U_I34051 ( .A(g25204), .ZN(I34051) );
INV_X32 U_g26159 ( .A(I34051), .ZN(g26159) );
INV_X32 U_I34056 ( .A(g25206), .ZN(I34056) );
INV_X32 U_g26164 ( .A(I34056), .ZN(g26164) );
INV_X32 U_I34059 ( .A(g25207), .ZN(I34059) );
INV_X32 U_g26165 ( .A(I34059), .ZN(g26165) );
INV_X32 U_I34063 ( .A(g25209), .ZN(I34063) );
INV_X32 U_g26167 ( .A(I34063), .ZN(g26167) );
INV_X32 U_I34068 ( .A(g25211), .ZN(I34068) );
INV_X32 U_g26172 ( .A(I34068), .ZN(g26172) );
INV_X32 U_I34071 ( .A(g25212), .ZN(I34071) );
INV_X32 U_g26173 ( .A(I34071), .ZN(g26173) );
INV_X32 U_I34074 ( .A(g25213), .ZN(I34074) );
INV_X32 U_g26174 ( .A(I34074), .ZN(g26174) );
INV_X32 U_I34077 ( .A(g25954), .ZN(I34077) );
INV_X32 U_g26175 ( .A(I34077), .ZN(g26175) );
INV_X32 U_I34080 ( .A(g25539), .ZN(I34080) );
INV_X32 U_g26178 ( .A(I34080), .ZN(g26178) );
INV_X32 U_I34083 ( .A(g25214), .ZN(I34083) );
INV_X32 U_g26181 ( .A(I34083), .ZN(g26181) );
INV_X32 U_I34086 ( .A(g25215), .ZN(I34086) );
INV_X32 U_g26182 ( .A(I34086), .ZN(g26182) );
INV_X32 U_I34091 ( .A(g25217), .ZN(I34091) );
INV_X32 U_g26187 ( .A(I34091), .ZN(g26187) );
INV_X32 U_g26189 ( .A(g25952), .ZN(g26189) );
INV_X32 U_I34096 ( .A(g25218), .ZN(I34096) );
INV_X32 U_g26190 ( .A(I34096), .ZN(g26190) );
INV_X32 U_I34099 ( .A(g25219), .ZN(I34099) );
INV_X32 U_g26191 ( .A(I34099), .ZN(g26191) );
INV_X32 U_I34102 ( .A(g25220), .ZN(I34102) );
INV_X32 U_g26192 ( .A(I34102), .ZN(g26192) );
INV_X32 U_I34105 ( .A(g25221), .ZN(I34105) );
INV_X32 U_g26193 ( .A(I34105), .ZN(g26193) );
INV_X32 U_I34108 ( .A(g25222), .ZN(I34108) );
INV_X32 U_g26194 ( .A(I34108), .ZN(g26194) );
INV_X32 U_I34111 ( .A(g25223), .ZN(I34111) );
INV_X32 U_g26195 ( .A(I34111), .ZN(g26195) );
INV_X32 U_I34114 ( .A(g25958), .ZN(I34114) );
INV_X32 U_g26196 ( .A(I34114), .ZN(g26196) );
INV_X32 U_I34118 ( .A(g25605), .ZN(I34118) );
INV_X32 U_g26202 ( .A(I34118), .ZN(g26202) );
INV_X32 U_I34121 ( .A(g25224), .ZN(I34121) );
INV_X32 U_g26205 ( .A(I34121), .ZN(g26205) );
INV_X32 U_I34124 ( .A(g25225), .ZN(I34124) );
INV_X32 U_g26206 ( .A(I34124), .ZN(g26206) );
INV_X32 U_I34128 ( .A(g25227), .ZN(I34128) );
INV_X32 U_g26208 ( .A(I34128), .ZN(g26208) );
INV_X32 U_g26209 ( .A(g25296), .ZN(g26209) );
INV_X32 U_I34132 ( .A(g25228), .ZN(I34132) );
INV_X32 U_g26210 ( .A(I34132), .ZN(g26210) );
INV_X32 U_I34135 ( .A(g25229), .ZN(I34135) );
INV_X32 U_g26211 ( .A(I34135), .ZN(g26211) );
INV_X32 U_I34140 ( .A(g25230), .ZN(I34140) );
INV_X32 U_g26214 ( .A(I34140), .ZN(g26214) );
INV_X32 U_I34143 ( .A(g25231), .ZN(I34143) );
INV_X32 U_g26215 ( .A(I34143), .ZN(g26215) );
INV_X32 U_I34146 ( .A(g25232), .ZN(I34146) );
INV_X32 U_g26216 ( .A(I34146), .ZN(g26216) );
INV_X32 U_I34150 ( .A(g25233), .ZN(I34150) );
INV_X32 U_g26220 ( .A(I34150), .ZN(g26220) );
INV_X32 U_I34153 ( .A(g25234), .ZN(I34153) );
INV_X32 U_g26221 ( .A(I34153), .ZN(g26221) );
INV_X32 U_I34156 ( .A(g25235), .ZN(I34156) );
INV_X32 U_g26222 ( .A(I34156), .ZN(g26222) );
INV_X32 U_I34159 ( .A(g25964), .ZN(I34159) );
INV_X32 U_g26223 ( .A(I34159), .ZN(g26223) );
INV_X32 U_I34162 ( .A(g25684), .ZN(I34162) );
INV_X32 U_g26226 ( .A(I34162), .ZN(g26226) );
INV_X32 U_I34165 ( .A(g25236), .ZN(I34165) );
INV_X32 U_g26229 ( .A(I34165), .ZN(g26229) );
INV_X32 U_I34168 ( .A(g25237), .ZN(I34168) );
INV_X32 U_g26230 ( .A(I34168), .ZN(g26230) );
INV_X32 U_I34172 ( .A(g25239), .ZN(I34172) );
INV_X32 U_g26232 ( .A(I34172), .ZN(g26232) );
INV_X32 U_g26237 ( .A(g25306), .ZN(g26237) );
INV_X32 U_I34180 ( .A(g25240), .ZN(I34180) );
INV_X32 U_g26238 ( .A(I34180), .ZN(g26238) );
INV_X32 U_I34183 ( .A(g25241), .ZN(I34183) );
INV_X32 U_g26239 ( .A(I34183), .ZN(g26239) );
INV_X32 U_I34189 ( .A(g25242), .ZN(I34189) );
INV_X32 U_g26245 ( .A(I34189), .ZN(g26245) );
INV_X32 U_I34192 ( .A(g25243), .ZN(I34192) );
INV_X32 U_g26246 ( .A(I34192), .ZN(g26246) );
INV_X32 U_I34195 ( .A(g25244), .ZN(I34195) );
INV_X32 U_g26247 ( .A(I34195), .ZN(g26247) );
INV_X32 U_I34198 ( .A(g25245), .ZN(I34198) );
INV_X32 U_g26248 ( .A(I34198), .ZN(g26248) );
INV_X32 U_I34201 ( .A(g25246), .ZN(I34201) );
INV_X32 U_g26249 ( .A(I34201), .ZN(g26249) );
INV_X32 U_I34204 ( .A(g25247), .ZN(I34204) );
INV_X32 U_g26250 ( .A(I34204), .ZN(g26250) );
INV_X32 U_I34207 ( .A(g25969), .ZN(I34207) );
INV_X32 U_g26251 ( .A(I34207), .ZN(g26251) );
INV_X32 U_I34210 ( .A(g25761), .ZN(I34210) );
INV_X32 U_g26254 ( .A(I34210), .ZN(g26254) );
INV_X32 U_I34220 ( .A(g25248), .ZN(I34220) );
INV_X32 U_g26264 ( .A(I34220), .ZN(g26264) );
INV_X32 U_g26275 ( .A(g25315), .ZN(g26275) );
INV_X32 U_I34230 ( .A(g25249), .ZN(I34230) );
INV_X32 U_g26276 ( .A(I34230), .ZN(g26276) );
INV_X32 U_I34233 ( .A(g25250), .ZN(I34233) );
INV_X32 U_g26277 ( .A(I34233), .ZN(g26277) );
INV_X32 U_I34238 ( .A(g25251), .ZN(I34238) );
INV_X32 U_g26280 ( .A(I34238), .ZN(g26280) );
INV_X32 U_I34241 ( .A(g25252), .ZN(I34241) );
INV_X32 U_g26281 ( .A(I34241), .ZN(g26281) );
INV_X32 U_I34244 ( .A(g25253), .ZN(I34244) );
INV_X32 U_g26282 ( .A(I34244), .ZN(g26282) );
INV_X32 U_I34254 ( .A(g25185), .ZN(I34254) );
INV_X32 U_g26294 ( .A(I34254), .ZN(g26294) );
INV_X32 U_I34266 ( .A(g25255), .ZN(I34266) );
INV_X32 U_g26308 ( .A(I34266), .ZN(g26308) );
INV_X32 U_g26313 ( .A(g25324), .ZN(g26313) );
INV_X32 U_I34274 ( .A(g25256), .ZN(I34274) );
INV_X32 U_g26314 ( .A(I34274), .ZN(g26314) );
INV_X32 U_I34277 ( .A(g25257), .ZN(I34277) );
INV_X32 U_g26315 ( .A(I34277), .ZN(g26315) );
INV_X32 U_I34296 ( .A(g25189), .ZN(I34296) );
INV_X32 U_g26341 ( .A(I34296), .ZN(g26341) );
INV_X32 U_I34306 ( .A(g25259), .ZN(I34306) );
INV_X32 U_g26349 ( .A(I34306), .ZN(g26349) );
INV_X32 U_I34313 ( .A(g25265), .ZN(I34313) );
INV_X32 U_g26354 ( .A(I34313), .ZN(g26354) );
INV_X32 U_I34316 ( .A(g25191), .ZN(I34316) );
INV_X32 U_g26355 ( .A(I34316), .ZN(g26355) );
INV_X32 U_I34321 ( .A(g25928), .ZN(I34321) );
INV_X32 U_g26358 ( .A(I34321), .ZN(g26358) );
INV_X32 U_I34327 ( .A(g25260), .ZN(I34327) );
INV_X32 U_g26364 ( .A(I34327), .ZN(g26364) );
INV_X32 U_I34343 ( .A(g25194), .ZN(I34343) );
INV_X32 U_g26385 ( .A(I34343), .ZN(g26385) );
INV_X32 U_I34353 ( .A(g25927), .ZN(I34353) );
INV_X32 U_g26393 ( .A(I34353), .ZN(g26393) );
INV_X32 U_I34358 ( .A(g25262), .ZN(I34358) );
INV_X32 U_g26398 ( .A(I34358), .ZN(g26398) );
INV_X32 U_I34363 ( .A(g25930), .ZN(I34363) );
INV_X32 U_g26401 ( .A(I34363), .ZN(g26401) );
INV_X32 U_I34369 ( .A(g25263), .ZN(I34369) );
INV_X32 U_g26407 ( .A(I34369), .ZN(g26407) );
INV_X32 U_I34385 ( .A(g25197), .ZN(I34385) );
INV_X32 U_g26428 ( .A(I34385), .ZN(g26428) );
INV_X32 U_I34388 ( .A(g25200), .ZN(I34388) );
INV_X32 U_g26429 ( .A(I34388), .ZN(g26429) );
INV_X32 U_I34392 ( .A(g25266), .ZN(I34392) );
INV_X32 U_g26433 ( .A(I34392), .ZN(g26433) );
INV_X32 U_I34395 ( .A(g25929), .ZN(I34395) );
INV_X32 U_g26434 ( .A(I34395), .ZN(g26434) );
INV_X32 U_I34400 ( .A(g25267), .ZN(I34400) );
INV_X32 U_g26439 ( .A(I34400), .ZN(g26439) );
INV_X32 U_I34405 ( .A(g25933), .ZN(I34405) );
INV_X32 U_g26442 ( .A(I34405), .ZN(g26442) );
INV_X32 U_I34411 ( .A(g25268), .ZN(I34411) );
INV_X32 U_g26448 ( .A(I34411), .ZN(g26448) );
INV_X32 U_I34421 ( .A(g25203), .ZN(I34421) );
INV_X32 U_g26461 ( .A(I34421), .ZN(g26461) );
INV_X32 U_I34425 ( .A(g25270), .ZN(I34425) );
INV_X32 U_g26465 ( .A(I34425), .ZN(g26465) );
INV_X32 U_I34428 ( .A(g25931), .ZN(I34428) );
INV_X32 U_g26466 ( .A(I34428), .ZN(g26466) );
INV_X32 U_I34433 ( .A(g25271), .ZN(I34433) );
INV_X32 U_g26471 ( .A(I34433), .ZN(g26471) );
INV_X32 U_I34438 ( .A(g25936), .ZN(I34438) );
INV_X32 U_g26474 ( .A(I34438), .ZN(g26474) );
INV_X32 U_I34444 ( .A(g25272), .ZN(I34444) );
INV_X32 U_g26480 ( .A(I34444), .ZN(g26480) );
INV_X32 U_g26481 ( .A(g25764), .ZN(g26481) );
INV_X32 U_I34449 ( .A(g25205), .ZN(I34449) );
INV_X32 U_g26485 ( .A(I34449), .ZN(g26485) );
INV_X32 U_I34453 ( .A(g25279), .ZN(I34453) );
INV_X32 U_g26489 ( .A(I34453), .ZN(g26489) );
INV_X32 U_I34456 ( .A(g25934), .ZN(I34456) );
INV_X32 U_g26490 ( .A(I34456), .ZN(g26490) );
INV_X32 U_I34461 ( .A(g25280), .ZN(I34461) );
INV_X32 U_g26495 ( .A(I34461), .ZN(g26495) );
INV_X32 U_I34464 ( .A(g25199), .ZN(I34464) );
INV_X32 U_g26496 ( .A(I34464), .ZN(g26496) );
INV_X32 U_g26497 ( .A(g25818), .ZN(g26497) );
INV_X32 U_I34469 ( .A(g25210), .ZN(I34469) );
INV_X32 U_g26501 ( .A(I34469), .ZN(g26501) );
INV_X32 U_I34473 ( .A(g25288), .ZN(I34473) );
INV_X32 U_g26505 ( .A(I34473), .ZN(g26505) );
INV_X32 U_I34476 ( .A(g25201), .ZN(I34476) );
INV_X32 U_g26506 ( .A(I34476), .ZN(g26506) );
INV_X32 U_I34479 ( .A(g25202), .ZN(I34479) );
INV_X32 U_g26507 ( .A(I34479), .ZN(g26507) );
INV_X32 U_g26508 ( .A(g25312), .ZN(g26508) );
INV_X32 U_g26512 ( .A(g25853), .ZN(g26512) );
INV_X32 U_g26516 ( .A(g25320), .ZN(g26516) );
INV_X32 U_g26520 ( .A(g25874), .ZN(g26520) );
INV_X32 U_g26521 ( .A(g25331), .ZN(g26521) );
INV_X32 U_g26525 ( .A(g25340), .ZN(g26525) );
INV_X32 U_g26533 ( .A(g25454), .ZN(g26533) );
INV_X32 U_g26538 ( .A(g25458), .ZN(g26538) );
INV_X32 U_g26539 ( .A(g25463), .ZN(g26539) );
INV_X32 U_g26540 ( .A(g25467), .ZN(g26540) );
INV_X32 U_g26542 ( .A(g25472), .ZN(g26542) );
INV_X32 U_g26543 ( .A(g25476), .ZN(g26543) );
INV_X32 U_g26544 ( .A(g25479), .ZN(g26544) );
INV_X32 U_g26546 ( .A(g25484), .ZN(g26546) );
INV_X32 U_I34505 ( .A(g25450), .ZN(I34505) );
INV_X32 U_g26548 ( .A(I34505), .ZN(g26548) );
INV_X32 U_g26549 ( .A(g25421), .ZN(g26549) );
INV_X32 U_g26550 ( .A(g25493), .ZN(g26550) );
INV_X32 U_g26551 ( .A(g25496), .ZN(g26551) );
INV_X32 U_g26552 ( .A(g25499), .ZN(g26552) );
INV_X32 U_g26554 ( .A(g25502), .ZN(g26554) );
INV_X32 U_g26555 ( .A(g25507), .ZN(g26555) );
INV_X32 U_g26556 ( .A(g25510), .ZN(g26556) );
INV_X32 U_g26558 ( .A(g25515), .ZN(g26558) );
INV_X32 U_g26561 ( .A(g25524), .ZN(g26561) );
INV_X32 U_g26562 ( .A(g25527), .ZN(g26562) );
INV_X32 U_g26563 ( .A(g25530), .ZN(g26563) );
INV_X32 U_g26564 ( .A(g25533), .ZN(g26564) );
INV_X32 U_g26565 ( .A(g25536), .ZN(g26565) );
INV_X32 U_g26566 ( .A(g25540), .ZN(g26566) );
INV_X32 U_g26567 ( .A(g25543), .ZN(g26567) );
INV_X32 U_g26568 ( .A(g25546), .ZN(g26568) );
INV_X32 U_g26570 ( .A(g25549), .ZN(g26570) );
INV_X32 U_g26571 ( .A(g25554), .ZN(g26571) );
INV_X32 U_g26572 ( .A(g25557), .ZN(g26572) );
INV_X32 U_g26574 ( .A(g25562), .ZN(g26574) );
INV_X32 U_I34535 ( .A(g25451), .ZN(I34535) );
INV_X32 U_g26576 ( .A(I34535), .ZN(g26576) );
INV_X32 U_g26577 ( .A(g25436), .ZN(g26577) );
INV_X32 U_g26578 ( .A(g25573), .ZN(g26578) );
INV_X32 U_g26579 ( .A(g25576), .ZN(g26579) );
INV_X32 U_g26580 ( .A(g25579), .ZN(g26580) );
INV_X32 U_g26581 ( .A(g25582), .ZN(g26581) );
INV_X32 U_g26582 ( .A(g25585), .ZN(g26582) );
INV_X32 U_g26584 ( .A(g25590), .ZN(g26584) );
INV_X32 U_g26585 ( .A(g25593), .ZN(g26585) );
INV_X32 U_g26586 ( .A(g25596), .ZN(g26586) );
INV_X32 U_g26587 ( .A(g25599), .ZN(g26587) );
INV_X32 U_g26588 ( .A(g25602), .ZN(g26588) );
INV_X32 U_g26589 ( .A(g25606), .ZN(g26589) );
INV_X32 U_g26590 ( .A(g25609), .ZN(g26590) );
INV_X32 U_g26591 ( .A(g25612), .ZN(g26591) );
INV_X32 U_g26593 ( .A(g25615), .ZN(g26593) );
INV_X32 U_g26594 ( .A(g25620), .ZN(g26594) );
INV_X32 U_g26595 ( .A(g25623), .ZN(g26595) );
INV_X32 U_g26597 ( .A(g25443), .ZN(g26597) );
INV_X32 U_g26598 ( .A(g25634), .ZN(g26598) );
INV_X32 U_g26599 ( .A(g25637), .ZN(g26599) );
INV_X32 U_g26600 ( .A(g25640), .ZN(g26600) );
INV_X32 U_g26601 ( .A(g25643), .ZN(g26601) );
INV_X32 U_g26602 ( .A(g25652), .ZN(g26602) );
INV_X32 U_g26603 ( .A(g25655), .ZN(g26603) );
INV_X32 U_g26604 ( .A(g25658), .ZN(g26604) );
INV_X32 U_g26605 ( .A(g25661), .ZN(g26605) );
INV_X32 U_g26606 ( .A(g25664), .ZN(g26606) );
INV_X32 U_g26608 ( .A(g25669), .ZN(g26608) );
INV_X32 U_g26609 ( .A(g25672), .ZN(g26609) );
INV_X32 U_g26610 ( .A(g25675), .ZN(g26610) );
INV_X32 U_g26611 ( .A(g25678), .ZN(g26611) );
INV_X32 U_g26612 ( .A(g25681), .ZN(g26612) );
INV_X32 U_g26613 ( .A(g25685), .ZN(g26613) );
INV_X32 U_g26614 ( .A(g25688), .ZN(g26614) );
INV_X32 U_g26615 ( .A(g25691), .ZN(g26615) );
INV_X32 U_g26617 ( .A(g25694), .ZN(g26617) );
INV_X32 U_I34579 ( .A(g25452), .ZN(I34579) );
INV_X32 U_g26618 ( .A(I34579), .ZN(g26618) );
INV_X32 U_g26619 ( .A(g25700), .ZN(g26619) );
INV_X32 U_g26620 ( .A(g25703), .ZN(g26620) );
INV_X32 U_g26621 ( .A(g25711), .ZN(g26621) );
INV_X32 U_g26622 ( .A(g25714), .ZN(g26622) );
INV_X32 U_g26623 ( .A(g25717), .ZN(g26623) );
INV_X32 U_g26624 ( .A(g25720), .ZN(g26624) );
INV_X32 U_g26625 ( .A(g25729), .ZN(g26625) );
INV_X32 U_g26626 ( .A(g25732), .ZN(g26626) );
INV_X32 U_g26627 ( .A(g25735), .ZN(g26627) );
INV_X32 U_g26628 ( .A(g25738), .ZN(g26628) );
INV_X32 U_g26629 ( .A(g25741), .ZN(g26629) );
INV_X32 U_g26631 ( .A(g25746), .ZN(g26631) );
INV_X32 U_g26632 ( .A(g25749), .ZN(g26632) );
INV_X32 U_g26633 ( .A(g25752), .ZN(g26633) );
INV_X32 U_g26634 ( .A(g25755), .ZN(g26634) );
INV_X32 U_g26635 ( .A(g25758), .ZN(g26635) );
INV_X32 U_g26636 ( .A(g25767), .ZN(g26636) );
INV_X32 U_g26637 ( .A(g25773), .ZN(g26637) );
INV_X32 U_g26638 ( .A(g25776), .ZN(g26638) );
INV_X32 U_g26639 ( .A(g25784), .ZN(g26639) );
INV_X32 U_g26640 ( .A(g25787), .ZN(g26640) );
INV_X32 U_g26641 ( .A(g25790), .ZN(g26641) );
INV_X32 U_g26642 ( .A(g25793), .ZN(g26642) );
INV_X32 U_g26643 ( .A(g25802), .ZN(g26643) );
INV_X32 U_g26644 ( .A(g25805), .ZN(g26644) );
INV_X32 U_g26645 ( .A(g25808), .ZN(g26645) );
INV_X32 U_g26646 ( .A(g25811), .ZN(g26646) );
INV_X32 U_g26647 ( .A(g25814), .ZN(g26647) );
INV_X32 U_g26648 ( .A(g25821), .ZN(g26648) );
INV_X32 U_g26649 ( .A(g25827), .ZN(g26649) );
INV_X32 U_g26650 ( .A(g25830), .ZN(g26650) );
INV_X32 U_g26651 ( .A(g25838), .ZN(g26651) );
INV_X32 U_g26652 ( .A(g25841), .ZN(g26652) );
INV_X32 U_g26653 ( .A(g25844), .ZN(g26653) );
INV_X32 U_g26654 ( .A(g25847), .ZN(g26654) );
INV_X32 U_g26656 ( .A(g25856), .ZN(g26656) );
INV_X32 U_g26657 ( .A(g25862), .ZN(g26657) );
INV_X32 U_g26658 ( .A(g25865), .ZN(g26658) );
INV_X32 U_g26662 ( .A(g25877), .ZN(g26662) );
INV_X32 U_I34641 ( .A(g26086), .ZN(I34641) );
INV_X32 U_g26678 ( .A(I34641), .ZN(g26678) );
INV_X32 U_I34644 ( .A(g26159), .ZN(I34644) );
INV_X32 U_g26679 ( .A(I34644), .ZN(g26679) );
INV_X32 U_I34647 ( .A(g26164), .ZN(I34647) );
INV_X32 U_g26680 ( .A(I34647), .ZN(g26680) );
INV_X32 U_I34650 ( .A(g26172), .ZN(I34650) );
INV_X32 U_g26681 ( .A(I34650), .ZN(g26681) );
INV_X32 U_I34653 ( .A(g26165), .ZN(I34653) );
INV_X32 U_g26682 ( .A(I34653), .ZN(g26682) );
INV_X32 U_I34656 ( .A(g26173), .ZN(I34656) );
INV_X32 U_g26683 ( .A(I34656), .ZN(g26683) );
INV_X32 U_I34659 ( .A(g26190), .ZN(I34659) );
INV_X32 U_g26684 ( .A(I34659), .ZN(g26684) );
INV_X32 U_I34662 ( .A(g26174), .ZN(I34662) );
INV_X32 U_g26685 ( .A(I34662), .ZN(g26685) );
INV_X32 U_I34665 ( .A(g26191), .ZN(I34665) );
INV_X32 U_g26686 ( .A(I34665), .ZN(g26686) );
INV_X32 U_I34668 ( .A(g26210), .ZN(I34668) );
INV_X32 U_g26687 ( .A(I34668), .ZN(g26687) );
INV_X32 U_I34671 ( .A(g26192), .ZN(I34671) );
INV_X32 U_g26688 ( .A(I34671), .ZN(g26688) );
INV_X32 U_I34674 ( .A(g26211), .ZN(I34674) );
INV_X32 U_g26689 ( .A(I34674), .ZN(g26689) );
INV_X32 U_I34677 ( .A(g26232), .ZN(I34677) );
INV_X32 U_g26690 ( .A(I34677), .ZN(g26690) );
INV_X32 U_I34680 ( .A(g26294), .ZN(I34680) );
INV_X32 U_g26691 ( .A(I34680), .ZN(g26691) );
INV_X32 U_I34683 ( .A(g26364), .ZN(I34683) );
INV_X32 U_g26692 ( .A(I34683), .ZN(g26692) );
INV_X32 U_I34686 ( .A(g26398), .ZN(I34686) );
INV_X32 U_g26693 ( .A(I34686), .ZN(g26693) );
INV_X32 U_I34689 ( .A(g26433), .ZN(I34689) );
INV_X32 U_g26694 ( .A(I34689), .ZN(g26694) );
INV_X32 U_I34692 ( .A(g26102), .ZN(I34692) );
INV_X32 U_g26695 ( .A(I34692), .ZN(g26695) );
INV_X32 U_I34695 ( .A(g26167), .ZN(I34695) );
INV_X32 U_g26696 ( .A(I34695), .ZN(g26696) );
INV_X32 U_I34698 ( .A(g26181), .ZN(I34698) );
INV_X32 U_g26697 ( .A(I34698), .ZN(g26697) );
INV_X32 U_I34701 ( .A(g26193), .ZN(I34701) );
INV_X32 U_g26698 ( .A(I34701), .ZN(g26698) );
INV_X32 U_I34704 ( .A(g26182), .ZN(I34704) );
INV_X32 U_g26699 ( .A(I34704), .ZN(g26699) );
INV_X32 U_I34707 ( .A(g26194), .ZN(I34707) );
INV_X32 U_g26700 ( .A(I34707), .ZN(g26700) );
INV_X32 U_I34710 ( .A(g26214), .ZN(I34710) );
INV_X32 U_g26701 ( .A(I34710), .ZN(g26701) );
INV_X32 U_I34713 ( .A(g26195), .ZN(I34713) );
INV_X32 U_g26702 ( .A(I34713), .ZN(g26702) );
INV_X32 U_I34716 ( .A(g26215), .ZN(I34716) );
INV_X32 U_g26703 ( .A(I34716), .ZN(g26703) );
INV_X32 U_I34719 ( .A(g26238), .ZN(I34719) );
INV_X32 U_g26704 ( .A(I34719), .ZN(g26704) );
INV_X32 U_I34722 ( .A(g26216), .ZN(I34722) );
INV_X32 U_g26705 ( .A(I34722), .ZN(g26705) );
INV_X32 U_I34725 ( .A(g26239), .ZN(I34725) );
INV_X32 U_g26706 ( .A(I34725), .ZN(g26706) );
INV_X32 U_I34728 ( .A(g26264), .ZN(I34728) );
INV_X32 U_g26707 ( .A(I34728), .ZN(g26707) );
INV_X32 U_I34731 ( .A(g26341), .ZN(I34731) );
INV_X32 U_g26708 ( .A(I34731), .ZN(g26708) );
INV_X32 U_I34734 ( .A(g26407), .ZN(I34734) );
INV_X32 U_g26709 ( .A(I34734), .ZN(g26709) );
INV_X32 U_I34737 ( .A(g26439), .ZN(I34737) );
INV_X32 U_g26710 ( .A(I34737), .ZN(g26710) );
INV_X32 U_I34740 ( .A(g26465), .ZN(I34740) );
INV_X32 U_g26711 ( .A(I34740), .ZN(g26711) );
INV_X32 U_I34743 ( .A(g26118), .ZN(I34743) );
INV_X32 U_g26712 ( .A(I34743), .ZN(g26712) );
INV_X32 U_I34746 ( .A(g26187), .ZN(I34746) );
INV_X32 U_g26713 ( .A(I34746), .ZN(g26713) );
INV_X32 U_I34749 ( .A(g26205), .ZN(I34749) );
INV_X32 U_g26714 ( .A(I34749), .ZN(g26714) );
INV_X32 U_I34752 ( .A(g26220), .ZN(I34752) );
INV_X32 U_g26715 ( .A(I34752), .ZN(g26715) );
INV_X32 U_I34755 ( .A(g26206), .ZN(I34755) );
INV_X32 U_g26716 ( .A(I34755), .ZN(g26716) );
INV_X32 U_I34758 ( .A(g26221), .ZN(I34758) );
INV_X32 U_g26717 ( .A(I34758), .ZN(g26717) );
INV_X32 U_I34761 ( .A(g26245), .ZN(I34761) );
INV_X32 U_g26718 ( .A(I34761), .ZN(g26718) );
INV_X32 U_I34764 ( .A(g26222), .ZN(I34764) );
INV_X32 U_g26719 ( .A(I34764), .ZN(g26719) );
INV_X32 U_I34767 ( .A(g26246), .ZN(I34767) );
INV_X32 U_g26720 ( .A(I34767), .ZN(g26720) );
INV_X32 U_I34770 ( .A(g26276), .ZN(I34770) );
INV_X32 U_g26721 ( .A(I34770), .ZN(g26721) );
INV_X32 U_I34773 ( .A(g26247), .ZN(I34773) );
INV_X32 U_g26722 ( .A(I34773), .ZN(g26722) );
INV_X32 U_I34776 ( .A(g26277), .ZN(I34776) );
INV_X32 U_g26723 ( .A(I34776), .ZN(g26723) );
INV_X32 U_I34779 ( .A(g26308), .ZN(I34779) );
INV_X32 U_g26724 ( .A(I34779), .ZN(g26724) );
INV_X32 U_I34782 ( .A(g26385), .ZN(I34782) );
INV_X32 U_g26725 ( .A(I34782), .ZN(g26725) );
INV_X32 U_I34785 ( .A(g26448), .ZN(I34785) );
INV_X32 U_g26726 ( .A(I34785), .ZN(g26726) );
INV_X32 U_I34788 ( .A(g26471), .ZN(I34788) );
INV_X32 U_g26727 ( .A(I34788), .ZN(g26727) );
INV_X32 U_I34791 ( .A(g26489), .ZN(I34791) );
INV_X32 U_g26728 ( .A(I34791), .ZN(g26728) );
INV_X32 U_I34794 ( .A(g26125), .ZN(I34794) );
INV_X32 U_g26729 ( .A(I34794), .ZN(g26729) );
INV_X32 U_I34797 ( .A(g26208), .ZN(I34797) );
INV_X32 U_g26730 ( .A(I34797), .ZN(g26730) );
INV_X32 U_I34800 ( .A(g26229), .ZN(I34800) );
INV_X32 U_g26731 ( .A(I34800), .ZN(g26731) );
INV_X32 U_I34803 ( .A(g26248), .ZN(I34803) );
INV_X32 U_g26732 ( .A(I34803), .ZN(g26732) );
INV_X32 U_I34806 ( .A(g26230), .ZN(I34806) );
INV_X32 U_g26733 ( .A(I34806), .ZN(g26733) );
INV_X32 U_I34809 ( .A(g26249), .ZN(I34809) );
INV_X32 U_g26734 ( .A(I34809), .ZN(g26734) );
INV_X32 U_I34812 ( .A(g26280), .ZN(I34812) );
INV_X32 U_g26735 ( .A(I34812), .ZN(g26735) );
INV_X32 U_I34815 ( .A(g26250), .ZN(I34815) );
INV_X32 U_g26736 ( .A(I34815), .ZN(g26736) );
INV_X32 U_I34818 ( .A(g26281), .ZN(I34818) );
INV_X32 U_g26737 ( .A(I34818), .ZN(g26737) );
INV_X32 U_I34821 ( .A(g26314), .ZN(I34821) );
INV_X32 U_g26738 ( .A(I34821), .ZN(g26738) );
INV_X32 U_I34824 ( .A(g26282), .ZN(I34824) );
INV_X32 U_g26739 ( .A(I34824), .ZN(g26739) );
INV_X32 U_I34827 ( .A(g26315), .ZN(I34827) );
INV_X32 U_g26740 ( .A(I34827), .ZN(g26740) );
INV_X32 U_I34830 ( .A(g26349), .ZN(I34830) );
INV_X32 U_g26741 ( .A(I34830), .ZN(g26741) );
INV_X32 U_I34833 ( .A(g26428), .ZN(I34833) );
INV_X32 U_g26742 ( .A(I34833), .ZN(g26742) );
INV_X32 U_I34836 ( .A(g26480), .ZN(I34836) );
INV_X32 U_g26743 ( .A(I34836), .ZN(g26743) );
INV_X32 U_I34839 ( .A(g26495), .ZN(I34839) );
INV_X32 U_g26744 ( .A(I34839), .ZN(g26744) );
INV_X32 U_I34842 ( .A(g26505), .ZN(I34842) );
INV_X32 U_g26745 ( .A(I34842), .ZN(g26745) );
INV_X32 U_I34845 ( .A(g26496), .ZN(I34845) );
INV_X32 U_g26746 ( .A(I34845), .ZN(g26746) );
INV_X32 U_I34848 ( .A(g26506), .ZN(I34848) );
INV_X32 U_g26747 ( .A(I34848), .ZN(g26747) );
INV_X32 U_I34851 ( .A(g26354), .ZN(I34851) );
INV_X32 U_g26748 ( .A(I34851), .ZN(g26748) );
INV_X32 U_I34854 ( .A(g26507), .ZN(I34854) );
INV_X32 U_g26749 ( .A(I34854), .ZN(g26749) );
INV_X32 U_I34857 ( .A(g26355), .ZN(I34857) );
INV_X32 U_g26750 ( .A(I34857), .ZN(g26750) );
INV_X32 U_I34860 ( .A(g26548), .ZN(I34860) );
INV_X32 U_g26751 ( .A(I34860), .ZN(g26751) );
INV_X32 U_I34863 ( .A(g26576), .ZN(I34863) );
INV_X32 U_g26752 ( .A(I34863), .ZN(g26752) );
INV_X32 U_I34866 ( .A(g26618), .ZN(I34866) );
INV_X32 U_g26753 ( .A(I34866), .ZN(g26753) );
INV_X32 U_I34872 ( .A(g26217), .ZN(I34872) );
INV_X32 U_g26757 ( .A(I34872), .ZN(g26757) );
INV_X32 U_I34879 ( .A(g26240), .ZN(I34879) );
INV_X32 U_g26762 ( .A(I34879), .ZN(g26762) );
INV_X32 U_I34901 ( .A(g26295), .ZN(I34901) );
INV_X32 U_g26782 ( .A(I34901), .ZN(g26782) );
INV_X32 U_I34909 ( .A(g26265), .ZN(I34909) );
INV_X32 U_g26788 ( .A(I34909), .ZN(g26788) );
INV_X32 U_I34916 ( .A(g26240), .ZN(I34916) );
INV_X32 U_g26793 ( .A(I34916), .ZN(g26793) );
INV_X32 U_I34921 ( .A(g26217), .ZN(I34921) );
INV_X32 U_g26796 ( .A(I34921), .ZN(g26796) );
INV_X32 U_I34946 ( .A(g26534), .ZN(I34946) );
INV_X32 U_g26819 ( .A(I34946), .ZN(g26819) );
INV_X32 U_I34957 ( .A(g26541), .ZN(I34957) );
INV_X32 U_g26828 ( .A(I34957), .ZN(g26828) );
INV_X32 U_I34961 ( .A(g26545), .ZN(I34961) );
INV_X32 U_g26830 ( .A(I34961), .ZN(g26830) );
INV_X32 U_I34964 ( .A(g26547), .ZN(I34964) );
INV_X32 U_g26831 ( .A(I34964), .ZN(g26831) );
INV_X32 U_I34967 ( .A(g26553), .ZN(I34967) );
INV_X32 U_g26832 ( .A(I34967), .ZN(g26832) );
INV_X32 U_I34971 ( .A(g26557), .ZN(I34971) );
INV_X32 U_g26834 ( .A(I34971), .ZN(g26834) );
INV_X32 U_I34974 ( .A(g26168), .ZN(I34974) );
INV_X32 U_g26835 ( .A(I34974), .ZN(g26835) );
INV_X32 U_I34977 ( .A(g26559), .ZN(I34977) );
INV_X32 U_g26836 ( .A(I34977), .ZN(g26836) );
INV_X32 U_I34980 ( .A(g26458), .ZN(I34980) );
INV_X32 U_g26837 ( .A(I34980), .ZN(g26837) );
INV_X32 U_I34983 ( .A(g26569), .ZN(I34983) );
INV_X32 U_g26840 ( .A(I34983), .ZN(g26840) );
INV_X32 U_I34986 ( .A(g26160), .ZN(I34986) );
INV_X32 U_g26841 ( .A(I34986), .ZN(g26841) );
INV_X32 U_I34990 ( .A(g26573), .ZN(I34990) );
INV_X32 U_g26843 ( .A(I34990), .ZN(g26843) );
INV_X32 U_I34993 ( .A(g26575), .ZN(I34993) );
INV_X32 U_g26844 ( .A(I34993), .ZN(g26844) );
INV_X32 U_I34997 ( .A(g26482), .ZN(I34997) );
INV_X32 U_g26846 ( .A(I34997), .ZN(g26846) );
INV_X32 U_I35000 ( .A(g26336), .ZN(I35000) );
INV_X32 U_g26849 ( .A(I35000), .ZN(g26849) );
INV_X32 U_I35003 ( .A(g26592), .ZN(I35003) );
INV_X32 U_g26850 ( .A(I35003), .ZN(g26850) );
INV_X32 U_I35007 ( .A(g26596), .ZN(I35007) );
INV_X32 U_g26852 ( .A(I35007), .ZN(g26852) );
INV_X32 U_I35011 ( .A(g26304), .ZN(I35011) );
INV_X32 U_g26854 ( .A(I35011), .ZN(g26854) );
INV_X32 U_I35014 ( .A(g26498), .ZN(I35014) );
INV_X32 U_g26855 ( .A(I35014), .ZN(g26855) );
INV_X32 U_I35017 ( .A(g26616), .ZN(I35017) );
INV_X32 U_g26858 ( .A(I35017), .ZN(g26858) );
INV_X32 U_I35028 ( .A(g26513), .ZN(I35028) );
INV_X32 U_g26861 ( .A(I35028), .ZN(g26861) );
INV_X32 U_I35031 ( .A(g26529), .ZN(I35031) );
INV_X32 U_g26864 ( .A(I35031), .ZN(g26864) );
INV_X32 U_I35049 ( .A(g26530), .ZN(I35049) );
INV_X32 U_g26868 ( .A(I35049), .ZN(g26868) );
INV_X32 U_I35053 ( .A(g26655), .ZN(I35053) );
INV_X32 U_g26872 ( .A(I35053), .ZN(g26872) );
INV_X32 U_I35064 ( .A(g26531), .ZN(I35064) );
INV_X32 U_g26875 ( .A(I35064), .ZN(g26875) );
INV_X32 U_I35067 ( .A(g26659), .ZN(I35067) );
INV_X32 U_g26876 ( .A(I35067), .ZN(g26876) );
INV_X32 U_I35072 ( .A(g26661), .ZN(I35072) );
INV_X32 U_g26881 ( .A(I35072), .ZN(g26881) );
INV_X32 U_I35076 ( .A(g26532), .ZN(I35076) );
INV_X32 U_g26883 ( .A(I35076), .ZN(g26883) );
INV_X32 U_I35079 ( .A(g26664), .ZN(I35079) );
INV_X32 U_g26884 ( .A(I35079), .ZN(g26884) );
INV_X32 U_I35083 ( .A(g26665), .ZN(I35083) );
INV_X32 U_g26886 ( .A(I35083), .ZN(g26886) );
INV_X32 U_I35087 ( .A(g26667), .ZN(I35087) );
INV_X32 U_g26890 ( .A(I35087), .ZN(g26890) );
INV_X32 U_I35092 ( .A(g26669), .ZN(I35092) );
INV_X32 U_g26895 ( .A(I35092), .ZN(g26895) );
INV_X32 U_I35095 ( .A(g26670), .ZN(I35095) );
INV_X32 U_g26896 ( .A(I35095), .ZN(g26896) );
INV_X32 U_I35099 ( .A(g26672), .ZN(I35099) );
INV_X32 U_g26900 ( .A(I35099), .ZN(g26900) );
INV_X32 U_I35106 ( .A(g26675), .ZN(I35106) );
INV_X32 U_g26909 ( .A(I35106), .ZN(g26909) );
INV_X32 U_I35109 ( .A(g26676), .ZN(I35109) );
INV_X32 U_g26910 ( .A(I35109), .ZN(g26910) );
INV_X32 U_I35116 ( .A(g26025), .ZN(I35116) );
INV_X32 U_g26921 ( .A(I35116), .ZN(g26921) );
INV_X32 U_g26922 ( .A(g26283), .ZN(g26922) );
INV_X32 U_g26935 ( .A(g26327), .ZN(g26935) );
INV_X32 U_g26944 ( .A(g26374), .ZN(g26944) );
INV_X32 U_g26950 ( .A(g26417), .ZN(g26950) );
INV_X32 U_I35136 ( .A(g26660), .ZN(I35136) );
INV_X32 U_g26953 ( .A(I35136), .ZN(g26953) );
INV_X32 U_g26954 ( .A(g26549), .ZN(g26954) );
INV_X32 U_I35141 ( .A(g26666), .ZN(I35141) );
INV_X32 U_g26956 ( .A(I35141), .ZN(g26956) );
INV_X32 U_g26957 ( .A(g26577), .ZN(g26957) );
INV_X32 U_I35146 ( .A(g26671), .ZN(I35146) );
INV_X32 U_g26959 ( .A(I35146), .ZN(g26959) );
INV_X32 U_g26960 ( .A(g26597), .ZN(g26960) );
INV_X32 U_I35153 ( .A(g26677), .ZN(I35153) );
INV_X32 U_g26964 ( .A(I35153), .ZN(g26964) );
INV_X32 U_I35172 ( .A(g26272), .ZN(I35172) );
INV_X32 U_g26983 ( .A(I35172), .ZN(g26983) );
INV_X32 U_g26987 ( .A(g26056), .ZN(g26987) );
INV_X32 U_g27010 ( .A(g26063), .ZN(g27010) );
INV_X32 U_g27036 ( .A(g26070), .ZN(g27036) );
INV_X32 U_g27064 ( .A(g26076), .ZN(g27064) );
INV_X32 U_I35254 ( .A(g26048), .ZN(I35254) );
INV_X32 U_g27075 ( .A(I35254), .ZN(g27075) );
INV_X32 U_I35283 ( .A(g26031), .ZN(I35283) );
INV_X32 U_g27102 ( .A(I35283), .ZN(g27102) );
INV_X32 U_I35297 ( .A(g26199), .ZN(I35297) );
INV_X32 U_g27114 ( .A(I35297), .ZN(g27114) );
INV_X32 U_I35301 ( .A(g26037), .ZN(I35301) );
INV_X32 U_g27116 ( .A(I35301), .ZN(g27116) );
INV_X32 U_I35313 ( .A(g26534), .ZN(I35313) );
INV_X32 U_g27126 ( .A(I35313), .ZN(g27126) );
INV_X32 U_I35319 ( .A(g26183), .ZN(I35319) );
INV_X32 U_g27132 ( .A(I35319), .ZN(g27132) );
INV_X32 U_g27133 ( .A(g26105), .ZN(g27133) );
INV_X32 U_g27134 ( .A(g26175), .ZN(g27134) );
INV_X32 U_g27135 ( .A(g26178), .ZN(g27135) );
INV_X32 U_g27136 ( .A(g26196), .ZN(g27136) );
INV_X32 U_g27137 ( .A(g26202), .ZN(g27137) );
INV_X32 U_g27138 ( .A(g26223), .ZN(g27138) );
INV_X32 U_g27139 ( .A(g26226), .ZN(g27139) );
INV_X32 U_g27140 ( .A(g26136), .ZN(g27140) );
INV_X32 U_g27141 ( .A(g26251), .ZN(g27141) );
INV_X32 U_g27142 ( .A(g26254), .ZN(g27142) );
INV_X32 U_g27143 ( .A(g26150), .ZN(g27143) );
INV_X32 U_I35334 ( .A(g26106), .ZN(I35334) );
INV_X32 U_g27145 ( .A(I35334), .ZN(g27145) );
INV_X32 U_g27146 ( .A(g26358), .ZN(g27146) );
INV_X32 U_g27148 ( .A(g26393), .ZN(g27148) );
INV_X32 U_I35341 ( .A(g26120), .ZN(I35341) );
INV_X32 U_g27150 ( .A(I35341), .ZN(g27150) );
INV_X32 U_g27151 ( .A(g26401), .ZN(g27151) );
INV_X32 U_g27153 ( .A(g26429), .ZN(g27153) );
INV_X32 U_I35347 ( .A(g26265), .ZN(I35347) );
INV_X32 U_g27154 ( .A(I35347), .ZN(g27154) );
INV_X32 U_g27155 ( .A(g26434), .ZN(g27155) );
INV_X32 U_I35351 ( .A(g26272), .ZN(I35351) );
INV_X32 U_g27156 ( .A(I35351), .ZN(g27156) );
INV_X32 U_I35355 ( .A(g26130), .ZN(I35355) );
INV_X32 U_g27158 ( .A(I35355), .ZN(g27158) );
INV_X32 U_g27159 ( .A(g26442), .ZN(g27159) );
INV_X32 U_I35360 ( .A(g26295), .ZN(I35360) );
INV_X32 U_g27161 ( .A(I35360), .ZN(g27161) );
INV_X32 U_g27162 ( .A(g26461), .ZN(g27162) );
INV_X32 U_I35364 ( .A(g26304), .ZN(I35364) );
INV_X32 U_g27163 ( .A(I35364), .ZN(g27163) );
INV_X32 U_g27164 ( .A(g26466), .ZN(g27164) );
INV_X32 U_I35369 ( .A(g26144), .ZN(I35369) );
INV_X32 U_g27166 ( .A(I35369), .ZN(g27166) );
INV_X32 U_g27167 ( .A(g26474), .ZN(g27167) );
INV_X32 U_I35373 ( .A(g26189), .ZN(I35373) );
INV_X32 U_g27168 ( .A(I35373), .ZN(g27168) );
INV_X32 U_I35376 ( .A(g26336), .ZN(I35376) );
INV_X32 U_g27171 ( .A(I35376), .ZN(g27171) );
INV_X32 U_g27172 ( .A(g26485), .ZN(g27172) );
INV_X32 U_g27173 ( .A(g26490), .ZN(g27173) );
INV_X32 U_I35383 ( .A(g26160), .ZN(I35383) );
INV_X32 U_g27176 ( .A(I35383), .ZN(g27176) );
INV_X32 U_g27177 ( .A(g26501), .ZN(g27177) );
INV_X32 U_I35389 ( .A(g26168), .ZN(I35389) );
INV_X32 U_g27180 ( .A(I35389), .ZN(g27180) );
INV_X32 U_I35394 ( .A(g26183), .ZN(I35394) );
INV_X32 U_g27183 ( .A(I35394), .ZN(g27183) );
INV_X32 U_I35399 ( .A(g26199), .ZN(I35399) );
INV_X32 U_g27186 ( .A(I35399), .ZN(g27186) );
INV_X32 U_I35404 ( .A(g26864), .ZN(I35404) );
INV_X32 U_g27189 ( .A(I35404), .ZN(g27189) );
INV_X32 U_I35407 ( .A(g27145), .ZN(I35407) );
INV_X32 U_g27190 ( .A(I35407), .ZN(g27190) );
INV_X32 U_I35410 ( .A(g26872), .ZN(I35410) );
INV_X32 U_g27191 ( .A(I35410), .ZN(g27191) );
INV_X32 U_I35413 ( .A(g26876), .ZN(I35413) );
INV_X32 U_g27192 ( .A(I35413), .ZN(g27192) );
INV_X32 U_I35416 ( .A(g26884), .ZN(I35416) );
INV_X32 U_g27193 ( .A(I35416), .ZN(g27193) );
INV_X32 U_I35419 ( .A(g26828), .ZN(I35419) );
INV_X32 U_g27194 ( .A(I35419), .ZN(g27194) );
INV_X32 U_I35422 ( .A(g26830), .ZN(I35422) );
INV_X32 U_g27195 ( .A(I35422), .ZN(g27195) );
INV_X32 U_I35425 ( .A(g26832), .ZN(I35425) );
INV_X32 U_g27196 ( .A(I35425), .ZN(g27196) );
INV_X32 U_I35428 ( .A(g26953), .ZN(I35428) );
INV_X32 U_g27197 ( .A(I35428), .ZN(g27197) );
INV_X32 U_I35431 ( .A(g26868), .ZN(I35431) );
INV_X32 U_g27198 ( .A(I35431), .ZN(g27198) );
INV_X32 U_I35434 ( .A(g27150), .ZN(I35434) );
INV_X32 U_g27199 ( .A(I35434), .ZN(g27199) );
INV_X32 U_I35437 ( .A(g27183), .ZN(I35437) );
INV_X32 U_g27200 ( .A(I35437), .ZN(g27200) );
INV_X32 U_I35440 ( .A(g27186), .ZN(I35440) );
INV_X32 U_g27201 ( .A(I35440), .ZN(g27201) );
INV_X32 U_I35443 ( .A(g26757), .ZN(I35443) );
INV_X32 U_g27202 ( .A(I35443), .ZN(g27202) );
INV_X32 U_I35446 ( .A(g26762), .ZN(I35446) );
INV_X32 U_g27203 ( .A(I35446), .ZN(g27203) );
INV_X32 U_I35449 ( .A(g27154), .ZN(I35449) );
INV_X32 U_g27204 ( .A(I35449), .ZN(g27204) );
INV_X32 U_I35452 ( .A(g27161), .ZN(I35452) );
INV_X32 U_g27205 ( .A(I35452), .ZN(g27205) );
INV_X32 U_I35455 ( .A(g26881), .ZN(I35455) );
INV_X32 U_g27206 ( .A(I35455), .ZN(g27206) );
INV_X32 U_I35458 ( .A(g26886), .ZN(I35458) );
INV_X32 U_g27207 ( .A(I35458), .ZN(g27207) );
INV_X32 U_I35461 ( .A(g26895), .ZN(I35461) );
INV_X32 U_g27208 ( .A(I35461), .ZN(g27208) );
INV_X32 U_I35464 ( .A(g26831), .ZN(I35464) );
INV_X32 U_g27209 ( .A(I35464), .ZN(g27209) );
INV_X32 U_I35467 ( .A(g26834), .ZN(I35467) );
INV_X32 U_g27210 ( .A(I35467), .ZN(g27210) );
INV_X32 U_I35470 ( .A(g26840), .ZN(I35470) );
INV_X32 U_g27211 ( .A(I35470), .ZN(g27211) );
INV_X32 U_I35473 ( .A(g27156), .ZN(I35473) );
INV_X32 U_g27212 ( .A(I35473), .ZN(g27212) );
INV_X32 U_I35476 ( .A(g27163), .ZN(I35476) );
INV_X32 U_g27213 ( .A(I35476), .ZN(g27213) );
INV_X32 U_I35479 ( .A(g27171), .ZN(I35479) );
INV_X32 U_g27214 ( .A(I35479), .ZN(g27214) );
INV_X32 U_I35482 ( .A(g27176), .ZN(I35482) );
INV_X32 U_g27215 ( .A(I35482), .ZN(g27215) );
INV_X32 U_I35485 ( .A(g27180), .ZN(I35485) );
INV_X32 U_g27216 ( .A(I35485), .ZN(g27216) );
INV_X32 U_I35488 ( .A(g26819), .ZN(I35488) );
INV_X32 U_g27217 ( .A(I35488), .ZN(g27217) );
INV_X32 U_I35491 ( .A(g26956), .ZN(I35491) );
INV_X32 U_g27218 ( .A(I35491), .ZN(g27218) );
INV_X32 U_I35494 ( .A(g26875), .ZN(I35494) );
INV_X32 U_g27219 ( .A(I35494), .ZN(g27219) );
INV_X32 U_I35497 ( .A(g27158), .ZN(I35497) );
INV_X32 U_g27220 ( .A(I35497), .ZN(g27220) );
INV_X32 U_I35500 ( .A(g26890), .ZN(I35500) );
INV_X32 U_g27221 ( .A(I35500), .ZN(g27221) );
INV_X32 U_I35503 ( .A(g26896), .ZN(I35503) );
INV_X32 U_g27222 ( .A(I35503), .ZN(g27222) );
INV_X32 U_I35506 ( .A(g26909), .ZN(I35506) );
INV_X32 U_g27223 ( .A(I35506), .ZN(g27223) );
INV_X32 U_I35509 ( .A(g26836), .ZN(I35509) );
INV_X32 U_g27224 ( .A(I35509), .ZN(g27224) );
INV_X32 U_I35512 ( .A(g26843), .ZN(I35512) );
INV_X32 U_g27225 ( .A(I35512), .ZN(g27225) );
INV_X32 U_I35515 ( .A(g26850), .ZN(I35515) );
INV_X32 U_g27226 ( .A(I35515), .ZN(g27226) );
INV_X32 U_I35518 ( .A(g26959), .ZN(I35518) );
INV_X32 U_g27227 ( .A(I35518), .ZN(g27227) );
INV_X32 U_I35521 ( .A(g26883), .ZN(I35521) );
INV_X32 U_g27228 ( .A(I35521), .ZN(g27228) );
INV_X32 U_I35524 ( .A(g27166), .ZN(I35524) );
INV_X32 U_g27229 ( .A(I35524), .ZN(g27229) );
INV_X32 U_I35527 ( .A(g26900), .ZN(I35527) );
INV_X32 U_g27230 ( .A(I35527), .ZN(g27230) );
INV_X32 U_I35530 ( .A(g26910), .ZN(I35530) );
INV_X32 U_g27231 ( .A(I35530), .ZN(g27231) );
INV_X32 U_I35533 ( .A(g26921), .ZN(I35533) );
INV_X32 U_g27232 ( .A(I35533), .ZN(g27232) );
INV_X32 U_I35536 ( .A(g26844), .ZN(I35536) );
INV_X32 U_g27233 ( .A(I35536), .ZN(g27233) );
INV_X32 U_I35539 ( .A(g26852), .ZN(I35539) );
INV_X32 U_g27234 ( .A(I35539), .ZN(g27234) );
INV_X32 U_I35542 ( .A(g26858), .ZN(I35542) );
INV_X32 U_g27235 ( .A(I35542), .ZN(g27235) );
INV_X32 U_I35545 ( .A(g26964), .ZN(I35545) );
INV_X32 U_g27236 ( .A(I35545), .ZN(g27236) );
INV_X32 U_I35548 ( .A(g27116), .ZN(I35548) );
INV_X32 U_g27237 ( .A(I35548), .ZN(g27237) );
INV_X32 U_I35551 ( .A(g27075), .ZN(I35551) );
INV_X32 U_g27238 ( .A(I35551), .ZN(g27238) );
INV_X32 U_I35554 ( .A(g27102), .ZN(I35554) );
INV_X32 U_g27239 ( .A(I35554), .ZN(g27239) );
INV_X32 U_g27349 ( .A(g27126), .ZN(g27349) );
INV_X32 U_I35667 ( .A(g27120), .ZN(I35667) );
INV_X32 U_g27353 ( .A(I35667), .ZN(g27353) );
INV_X32 U_I35673 ( .A(g27123), .ZN(I35673) );
INV_X32 U_g27357 ( .A(I35673), .ZN(g27357) );
INV_X32 U_I35678 ( .A(g27129), .ZN(I35678) );
INV_X32 U_g27360 ( .A(I35678), .ZN(g27360) );
INV_X32 U_I35681 ( .A(g26869), .ZN(I35681) );
INV_X32 U_g27361 ( .A(I35681), .ZN(g27361) );
INV_X32 U_I35686 ( .A(g27131), .ZN(I35686) );
INV_X32 U_g27366 ( .A(I35686), .ZN(g27366) );
INV_X32 U_I35689 ( .A(g26878), .ZN(I35689) );
INV_X32 U_g27367 ( .A(I35689), .ZN(g27367) );
INV_X32 U_I35695 ( .A(g26887), .ZN(I35695) );
INV_X32 U_g27373 ( .A(I35695), .ZN(g27373) );
INV_X32 U_I35698 ( .A(g26897), .ZN(I35698) );
INV_X32 U_g27376 ( .A(I35698), .ZN(g27376) );
INV_X32 U_I35708 ( .A(g26974), .ZN(I35708) );
INV_X32 U_g27380 ( .A(I35708), .ZN(g27380) );
INV_X32 U_I35711 ( .A(g26974), .ZN(I35711) );
INV_X32 U_g27381 ( .A(I35711), .ZN(g27381) );
INV_X32 U_g27383 ( .A(g27133), .ZN(g27383) );
INV_X32 U_g27384 ( .A(g27140), .ZN(g27384) );
INV_X32 U_I35723 ( .A(g27168), .ZN(I35723) );
INV_X32 U_g27385 ( .A(I35723), .ZN(g27385) );
INV_X32 U_g27386 ( .A(g27143), .ZN(g27386) );
INV_X32 U_I35727 ( .A(g26902), .ZN(I35727) );
INV_X32 U_g27387 ( .A(I35727), .ZN(g27387) );
INV_X32 U_I35731 ( .A(g26892), .ZN(I35731) );
INV_X32 U_g27391 ( .A(I35731), .ZN(g27391) );
INV_X32 U_I35737 ( .A(g26915), .ZN(I35737) );
INV_X32 U_g27397 ( .A(I35737), .ZN(g27397) );
INV_X32 U_I35741 ( .A(g27118), .ZN(I35741) );
INV_X32 U_g27401 ( .A(I35741), .ZN(g27401) );
INV_X32 U_I35744 ( .A(g26906), .ZN(I35744) );
INV_X32 U_g27404 ( .A(I35744), .ZN(g27404) );
INV_X32 U_I35750 ( .A(g26928), .ZN(I35750) );
INV_X32 U_g27410 ( .A(I35750), .ZN(g27410) );
INV_X32 U_I35756 ( .A(g27117), .ZN(I35756) );
INV_X32 U_g27416 ( .A(I35756), .ZN(g27416) );
INV_X32 U_I35759 ( .A(g27121), .ZN(I35759) );
INV_X32 U_g27419 ( .A(I35759), .ZN(g27419) );
INV_X32 U_I35762 ( .A(g26918), .ZN(I35762) );
INV_X32 U_g27422 ( .A(I35762), .ZN(g27422) );
INV_X32 U_I35768 ( .A(g26941), .ZN(I35768) );
INV_X32 U_g27428 ( .A(I35768), .ZN(g27428) );
INV_X32 U_I35772 ( .A(g26772), .ZN(I35772) );
INV_X32 U_g27432 ( .A(I35772), .ZN(g27432) );
INV_X32 U_I35777 ( .A(g27119), .ZN(I35777) );
INV_X32 U_g27437 ( .A(I35777), .ZN(g27437) );
INV_X32 U_I35780 ( .A(g27124), .ZN(I35780) );
INV_X32 U_g27440 ( .A(I35780), .ZN(g27440) );
INV_X32 U_I35783 ( .A(g26931), .ZN(I35783) );
INV_X32 U_g27443 ( .A(I35783), .ZN(g27443) );
INV_X32 U_g27449 ( .A(g26837), .ZN(g27449) );
INV_X32 U_I35791 ( .A(g26779), .ZN(I35791) );
INV_X32 U_g27451 ( .A(I35791), .ZN(g27451) );
INV_X32 U_I35796 ( .A(g27122), .ZN(I35796) );
INV_X32 U_g27456 ( .A(I35796), .ZN(g27456) );
INV_X32 U_I35799 ( .A(g27130), .ZN(I35799) );
INV_X32 U_g27459 ( .A(I35799), .ZN(g27459) );
INV_X32 U_I35803 ( .A(g26803), .ZN(I35803) );
INV_X32 U_g27463 ( .A(I35803), .ZN(g27463) );
INV_X32 U_g27465 ( .A(g26846), .ZN(g27465) );
INV_X32 U_I35809 ( .A(g26785), .ZN(I35809) );
INV_X32 U_g27467 ( .A(I35809), .ZN(g27467) );
INV_X32 U_I35814 ( .A(g27125), .ZN(I35814) );
INV_X32 U_g27472 ( .A(I35814), .ZN(g27472) );
INV_X32 U_I35817 ( .A(g26922), .ZN(I35817) );
INV_X32 U_g27475 ( .A(I35817), .ZN(g27475) );
INV_X32 U_I35821 ( .A(g26804), .ZN(I35821) );
INV_X32 U_g27479 ( .A(I35821), .ZN(g27479) );
INV_X32 U_I35824 ( .A(g26805), .ZN(I35824) );
INV_X32 U_g27480 ( .A(I35824), .ZN(g27480) );
INV_X32 U_I35829 ( .A(g26806), .ZN(I35829) );
INV_X32 U_g27483 ( .A(I35829), .ZN(g27483) );
INV_X32 U_g27484 ( .A(g26855), .ZN(g27484) );
INV_X32 U_I35834 ( .A(g26792), .ZN(I35834) );
INV_X32 U_g27486 ( .A(I35834), .ZN(g27486) );
INV_X32 U_I35837 ( .A(g26911), .ZN(I35837) );
INV_X32 U_g27489 ( .A(I35837), .ZN(g27489) );
INV_X32 U_I35841 ( .A(g26807), .ZN(I35841) );
INV_X32 U_g27493 ( .A(I35841), .ZN(g27493) );
INV_X32 U_I35844 ( .A(g26808), .ZN(I35844) );
INV_X32 U_g27494 ( .A(I35844), .ZN(g27494) );
INV_X32 U_I35849 ( .A(g26776), .ZN(I35849) );
INV_X32 U_g27497 ( .A(I35849), .ZN(g27497) );
INV_X32 U_I35852 ( .A(g26935), .ZN(I35852) );
INV_X32 U_g27498 ( .A(I35852), .ZN(g27498) );
INV_X32 U_I35856 ( .A(g26809), .ZN(I35856) );
INV_X32 U_g27502 ( .A(I35856), .ZN(g27502) );
INV_X32 U_I35859 ( .A(g26810), .ZN(I35859) );
INV_X32 U_g27503 ( .A(I35859), .ZN(g27503) );
INV_X32 U_I35863 ( .A(g26811), .ZN(I35863) );
INV_X32 U_g27505 ( .A(I35863), .ZN(g27505) );
INV_X32 U_g27506 ( .A(g26861), .ZN(g27506) );
INV_X32 U_I35868 ( .A(g26812), .ZN(I35868) );
INV_X32 U_g27508 ( .A(I35868), .ZN(g27508) );
INV_X32 U_I35872 ( .A(g26925), .ZN(I35872) );
INV_X32 U_g27510 ( .A(I35872), .ZN(g27510) );
INV_X32 U_I35876 ( .A(g26813), .ZN(I35876) );
INV_X32 U_g27514 ( .A(I35876), .ZN(g27514) );
INV_X32 U_I35879 ( .A(g26814), .ZN(I35879) );
INV_X32 U_g27515 ( .A(I35879), .ZN(g27515) );
INV_X32 U_I35883 ( .A(g26781), .ZN(I35883) );
INV_X32 U_g27517 ( .A(I35883), .ZN(g27517) );
INV_X32 U_I35886 ( .A(g26944), .ZN(I35886) );
INV_X32 U_g27518 ( .A(I35886), .ZN(g27518) );
INV_X32 U_I35890 ( .A(g26815), .ZN(I35890) );
INV_X32 U_g27522 ( .A(I35890), .ZN(g27522) );
INV_X32 U_I35893 ( .A(g26816), .ZN(I35893) );
INV_X32 U_g27523 ( .A(I35893), .ZN(g27523) );
INV_X32 U_I35897 ( .A(g26817), .ZN(I35897) );
INV_X32 U_g27525 ( .A(I35897), .ZN(g27525) );
INV_X32 U_I35900 ( .A(g26786), .ZN(I35900) );
INV_X32 U_g27526 ( .A(I35900), .ZN(g27526) );
INV_X32 U_I35915 ( .A(g26818), .ZN(I35915) );
INV_X32 U_g27533 ( .A(I35915), .ZN(g27533) );
INV_X32 U_I35919 ( .A(g26938), .ZN(I35919) );
INV_X32 U_g27535 ( .A(I35919), .ZN(g27535) );
INV_X32 U_I35923 ( .A(g26820), .ZN(I35923) );
INV_X32 U_g27539 ( .A(I35923), .ZN(g27539) );
INV_X32 U_I35926 ( .A(g26821), .ZN(I35926) );
INV_X32 U_g27540 ( .A(I35926), .ZN(g27540) );
INV_X32 U_I35930 ( .A(g26789), .ZN(I35930) );
INV_X32 U_g27542 ( .A(I35930), .ZN(g27542) );
INV_X32 U_I35933 ( .A(g26950), .ZN(I35933) );
INV_X32 U_g27543 ( .A(I35933), .ZN(g27543) );
INV_X32 U_I35937 ( .A(g26822), .ZN(I35937) );
INV_X32 U_g27547 ( .A(I35937), .ZN(g27547) );
INV_X32 U_I35940 ( .A(g26823), .ZN(I35940) );
INV_X32 U_g27548 ( .A(I35940), .ZN(g27548) );
INV_X32 U_I35953 ( .A(g26824), .ZN(I35953) );
INV_X32 U_g27553 ( .A(I35953), .ZN(g27553) );
INV_X32 U_I35957 ( .A(g26947), .ZN(I35957) );
INV_X32 U_g27555 ( .A(I35957), .ZN(g27555) );
INV_X32 U_I35961 ( .A(g26825), .ZN(I35961) );
INV_X32 U_g27559 ( .A(I35961), .ZN(g27559) );
INV_X32 U_I35964 ( .A(g26826), .ZN(I35964) );
INV_X32 U_g27560 ( .A(I35964), .ZN(g27560) );
INV_X32 U_I35968 ( .A(g26795), .ZN(I35968) );
INV_X32 U_g27562 ( .A(I35968), .ZN(g27562) );
INV_X32 U_I35983 ( .A(g26827), .ZN(I35983) );
INV_X32 U_g27569 ( .A(I35983), .ZN(g27569) );
INV_X32 U_I36008 ( .A(g26798), .ZN(I36008) );
INV_X32 U_g27586 ( .A(I36008), .ZN(g27586) );
INV_X32 U_g27589 ( .A(g27168), .ZN(g27589) );
INV_X32 U_g27590 ( .A(g27144), .ZN(g27590) );
INV_X32 U_g27595 ( .A(g27149), .ZN(g27595) );
INV_X32 U_g27599 ( .A(g27147), .ZN(g27599) );
INV_X32 U_g27604 ( .A(g27157), .ZN(g27604) );
INV_X32 U_g27608 ( .A(g27152), .ZN(g27608) );
INV_X32 U_g27613 ( .A(g27165), .ZN(g27613) );
INV_X32 U_g27617 ( .A(g27160), .ZN(g27617) );
INV_X32 U_g27622 ( .A(g27174), .ZN(g27622) );
INV_X32 U_I36032 ( .A(g27113), .ZN(I36032) );
INV_X32 U_g27632 ( .A(I36032), .ZN(g27632) );
INV_X32 U_I36042 ( .A(g26960), .ZN(I36042) );
INV_X32 U_g27662 ( .A(I36042), .ZN(g27662) );
INV_X32 U_I36046 ( .A(g26957), .ZN(I36046) );
INV_X32 U_g27667 ( .A(I36046), .ZN(g27667) );
INV_X32 U_I36052 ( .A(g26954), .ZN(I36052) );
INV_X32 U_g27674 ( .A(I36052), .ZN(g27674) );
INV_X32 U_I36060 ( .A(g27353), .ZN(I36060) );
INV_X32 U_g27683 ( .A(I36060), .ZN(g27683) );
INV_X32 U_I36063 ( .A(g27463), .ZN(I36063) );
INV_X32 U_g27684 ( .A(I36063), .ZN(g27684) );
INV_X32 U_I36066 ( .A(g27479), .ZN(I36066) );
INV_X32 U_g27685 ( .A(I36066), .ZN(g27685) );
INV_X32 U_I36069 ( .A(g27493), .ZN(I36069) );
INV_X32 U_g27686 ( .A(I36069), .ZN(g27686) );
INV_X32 U_I36072 ( .A(g27480), .ZN(I36072) );
INV_X32 U_g27687 ( .A(I36072), .ZN(g27687) );
INV_X32 U_I36075 ( .A(g27494), .ZN(I36075) );
INV_X32 U_g27688 ( .A(I36075), .ZN(g27688) );
INV_X32 U_I36078 ( .A(g27508), .ZN(I36078) );
INV_X32 U_g27689 ( .A(I36078), .ZN(g27689) );
INV_X32 U_I36081 ( .A(g27497), .ZN(I36081) );
INV_X32 U_g27690 ( .A(I36081), .ZN(g27690) );
INV_X32 U_I36084 ( .A(g27357), .ZN(I36084) );
INV_X32 U_g27691 ( .A(I36084), .ZN(g27691) );
INV_X32 U_I36087 ( .A(g27483), .ZN(I36087) );
INV_X32 U_g27692 ( .A(I36087), .ZN(g27692) );
INV_X32 U_I36090 ( .A(g27502), .ZN(I36090) );
INV_X32 U_g27693 ( .A(I36090), .ZN(g27693) );
INV_X32 U_I36093 ( .A(g27514), .ZN(I36093) );
INV_X32 U_g27694 ( .A(I36093), .ZN(g27694) );
INV_X32 U_I36096 ( .A(g27503), .ZN(I36096) );
INV_X32 U_g27695 ( .A(I36096), .ZN(g27695) );
INV_X32 U_I36099 ( .A(g27515), .ZN(I36099) );
INV_X32 U_g27696 ( .A(I36099), .ZN(g27696) );
INV_X32 U_I36102 ( .A(g27533), .ZN(I36102) );
INV_X32 U_g27697 ( .A(I36102), .ZN(g27697) );
INV_X32 U_I36105 ( .A(g27517), .ZN(I36105) );
INV_X32 U_g27698 ( .A(I36105), .ZN(g27698) );
INV_X32 U_I36108 ( .A(g27360), .ZN(I36108) );
INV_X32 U_g27699 ( .A(I36108), .ZN(g27699) );
INV_X32 U_I36111 ( .A(g27505), .ZN(I36111) );
INV_X32 U_g27700 ( .A(I36111), .ZN(g27700) );
INV_X32 U_I36114 ( .A(g27522), .ZN(I36114) );
INV_X32 U_g27701 ( .A(I36114), .ZN(g27701) );
INV_X32 U_I36117 ( .A(g27539), .ZN(I36117) );
INV_X32 U_g27702 ( .A(I36117), .ZN(g27702) );
INV_X32 U_I36120 ( .A(g27523), .ZN(I36120) );
INV_X32 U_g27703 ( .A(I36120), .ZN(g27703) );
INV_X32 U_I36123 ( .A(g27540), .ZN(I36123) );
INV_X32 U_g27704 ( .A(I36123), .ZN(g27704) );
INV_X32 U_I36126 ( .A(g27553), .ZN(I36126) );
INV_X32 U_g27705 ( .A(I36126), .ZN(g27705) );
INV_X32 U_I36129 ( .A(g27542), .ZN(I36129) );
INV_X32 U_g27706 ( .A(I36129), .ZN(g27706) );
INV_X32 U_I36132 ( .A(g27366), .ZN(I36132) );
INV_X32 U_g27707 ( .A(I36132), .ZN(g27707) );
INV_X32 U_I36135 ( .A(g27525), .ZN(I36135) );
INV_X32 U_g27708 ( .A(I36135), .ZN(g27708) );
INV_X32 U_I36138 ( .A(g27547), .ZN(I36138) );
INV_X32 U_g27709 ( .A(I36138), .ZN(g27709) );
INV_X32 U_I36141 ( .A(g27559), .ZN(I36141) );
INV_X32 U_g27710 ( .A(I36141), .ZN(g27710) );
INV_X32 U_I36144 ( .A(g27548), .ZN(I36144) );
INV_X32 U_g27711 ( .A(I36144), .ZN(g27711) );
INV_X32 U_I36147 ( .A(g27560), .ZN(I36147) );
INV_X32 U_g27712 ( .A(I36147), .ZN(g27712) );
INV_X32 U_I36150 ( .A(g27569), .ZN(I36150) );
INV_X32 U_g27713 ( .A(I36150), .ZN(g27713) );
INV_X32 U_I36153 ( .A(g27562), .ZN(I36153) );
INV_X32 U_g27714 ( .A(I36153), .ZN(g27714) );
INV_X32 U_I36156 ( .A(g27586), .ZN(I36156) );
INV_X32 U_g27715 ( .A(I36156), .ZN(g27715) );
INV_X32 U_I36159 ( .A(g27526), .ZN(I36159) );
INV_X32 U_g27716 ( .A(I36159), .ZN(g27716) );
INV_X32 U_I36162 ( .A(g27385), .ZN(I36162) );
INV_X32 U_g27717 ( .A(I36162), .ZN(g27717) );
INV_X32 U_g27748 ( .A(g27632), .ZN(g27748) );
INV_X32 U_I36213 ( .A(g27571), .ZN(I36213) );
INV_X32 U_g27776 ( .A(I36213), .ZN(g27776) );
INV_X32 U_I36217 ( .A(g27580), .ZN(I36217) );
INV_X32 U_g27780 ( .A(I36217), .ZN(g27780) );
INV_X32 U_I36221 ( .A(g27662), .ZN(I36221) );
INV_X32 U_g27784 ( .A(I36221), .ZN(g27784) );
INV_X32 U_I36224 ( .A(g27589), .ZN(I36224) );
INV_X32 U_g27785 ( .A(I36224), .ZN(g27785) );
INV_X32 U_I36227 ( .A(g27594), .ZN(I36227) );
INV_X32 U_g27786 ( .A(I36227), .ZN(g27786) );
INV_X32 U_I36230 ( .A(g27583), .ZN(I36230) );
INV_X32 U_g27787 ( .A(I36230), .ZN(g27787) );
INV_X32 U_I36234 ( .A(g27667), .ZN(I36234) );
INV_X32 U_g27791 ( .A(I36234), .ZN(g27791) );
INV_X32 U_I36237 ( .A(g27662), .ZN(I36237) );
INV_X32 U_g27792 ( .A(I36237), .ZN(g27792) );
INV_X32 U_I36240 ( .A(g27603), .ZN(I36240) );
INV_X32 U_g27793 ( .A(I36240), .ZN(g27793) );
INV_X32 U_I36243 ( .A(g27587), .ZN(I36243) );
INV_X32 U_g27794 ( .A(I36243), .ZN(g27794) );
INV_X32 U_I36246 ( .A(g27674), .ZN(I36246) );
INV_X32 U_g27797 ( .A(I36246), .ZN(g27797) );
INV_X32 U_I36250 ( .A(g27612), .ZN(I36250) );
INV_X32 U_g27799 ( .A(I36250), .ZN(g27799) );
INV_X32 U_I36253 ( .A(g27674), .ZN(I36253) );
INV_X32 U_g27800 ( .A(I36253), .ZN(g27800) );
INV_X32 U_I36264 ( .A(g27621), .ZN(I36264) );
INV_X32 U_g27805 ( .A(I36264), .ZN(g27805) );
INV_X32 U_I36267 ( .A(g27395), .ZN(I36267) );
INV_X32 U_g27806 ( .A(I36267), .ZN(g27806) );
INV_X32 U_I36280 ( .A(g27390), .ZN(I36280) );
INV_X32 U_g27817 ( .A(I36280), .ZN(g27817) );
INV_X32 U_I36283 ( .A(g27408), .ZN(I36283) );
INV_X32 U_g27820 ( .A(I36283), .ZN(g27820) );
INV_X32 U_I36296 ( .A(g27626), .ZN(I36296) );
INV_X32 U_g27831 ( .A(I36296), .ZN(g27831) );
INV_X32 U_I36307 ( .A(g27400), .ZN(I36307) );
INV_X32 U_g27839 ( .A(I36307), .ZN(g27839) );
INV_X32 U_I36311 ( .A(g27426), .ZN(I36311) );
INV_X32 U_g27843 ( .A(I36311), .ZN(g27843) );
INV_X32 U_I36321 ( .A(g27627), .ZN(I36321) );
INV_X32 U_g27847 ( .A(I36321), .ZN(g27847) );
INV_X32 U_I36327 ( .A(g27413), .ZN(I36327) );
INV_X32 U_g27858 ( .A(I36327), .ZN(g27858) );
INV_X32 U_I36330 ( .A(g27447), .ZN(I36330) );
INV_X32 U_g27861 ( .A(I36330), .ZN(g27861) );
INV_X32 U_I36337 ( .A(g27628), .ZN(I36337) );
INV_X32 U_g27872 ( .A(I36337), .ZN(g27872) );
INV_X32 U_I36341 ( .A(g27431), .ZN(I36341) );
INV_X32 U_g27879 ( .A(I36341), .ZN(g27879) );
INV_X32 U_I36347 ( .A(g27630), .ZN(I36347) );
INV_X32 U_g27889 ( .A(I36347), .ZN(g27889) );
INV_X32 U_I36354 ( .A(g27662), .ZN(I36354) );
INV_X32 U_g27903 ( .A(I36354), .ZN(g27903) );
INV_X32 U_I36358 ( .A(g27672), .ZN(I36358) );
INV_X32 U_g27905 ( .A(I36358), .ZN(g27905) );
INV_X32 U_I36362 ( .A(g27667), .ZN(I36362) );
INV_X32 U_g27907 ( .A(I36362), .ZN(g27907) );
INV_X32 U_I36367 ( .A(g27678), .ZN(I36367) );
INV_X32 U_g27910 ( .A(I36367), .ZN(g27910) );
INV_X32 U_I36371 ( .A(g27674), .ZN(I36371) );
INV_X32 U_g27912 ( .A(I36371), .ZN(g27912) );
INV_X32 U_I36379 ( .A(g27682), .ZN(I36379) );
INV_X32 U_g27918 ( .A(I36379), .ZN(g27918) );
INV_X32 U_I36382 ( .A(g27563), .ZN(I36382) );
INV_X32 U_g27919 ( .A(I36382), .ZN(g27919) );
INV_X32 U_I36390 ( .A(g27243), .ZN(I36390) );
INV_X32 U_g27927 ( .A(I36390), .ZN(g27927) );
INV_X32 U_I36393 ( .A(g27572), .ZN(I36393) );
INV_X32 U_g27928 ( .A(I36393), .ZN(g27928) );
INV_X32 U_I36397 ( .A(g27574), .ZN(I36397) );
INV_X32 U_g27932 ( .A(I36397), .ZN(g27932) );
INV_X32 U_I36404 ( .A(g27450), .ZN(I36404) );
INV_X32 U_g27939 ( .A(I36404), .ZN(g27939) );
INV_X32 U_I36407 ( .A(g27581), .ZN(I36407) );
INV_X32 U_g27942 ( .A(I36407), .ZN(g27942) );
INV_X32 U_I36411 ( .A(g27582), .ZN(I36411) );
INV_X32 U_g27946 ( .A(I36411), .ZN(g27946) );
INV_X32 U_I36417 ( .A(g27462), .ZN(I36417) );
INV_X32 U_g27952 ( .A(I36417), .ZN(g27952) );
INV_X32 U_I36420 ( .A(g27253), .ZN(I36420) );
INV_X32 U_g27955 ( .A(I36420), .ZN(g27955) );
INV_X32 U_I36423 ( .A(g27466), .ZN(I36423) );
INV_X32 U_g27956 ( .A(I36423), .ZN(g27956) );
INV_X32 U_I36426 ( .A(g27584), .ZN(I36426) );
INV_X32 U_g27959 ( .A(I36426), .ZN(g27959) );
INV_X32 U_I36432 ( .A(g27585), .ZN(I36432) );
INV_X32 U_g27965 ( .A(I36432), .ZN(g27965) );
INV_X32 U_g27969 ( .A(g27361), .ZN(g27969) );
INV_X32 U_I36438 ( .A(g27255), .ZN(I36438) );
INV_X32 U_g27971 ( .A(I36438), .ZN(g27971) );
INV_X32 U_I36441 ( .A(g27256), .ZN(I36441) );
INV_X32 U_g27972 ( .A(I36441), .ZN(g27972) );
INV_X32 U_I36444 ( .A(g27482), .ZN(I36444) );
INV_X32 U_g27973 ( .A(I36444), .ZN(g27973) );
INV_X32 U_I36447 ( .A(g27257), .ZN(I36447) );
INV_X32 U_g27976 ( .A(I36447), .ZN(g27976) );
INV_X32 U_I36450 ( .A(g27485), .ZN(I36450) );
INV_X32 U_g27977 ( .A(I36450), .ZN(g27977) );
INV_X32 U_I36454 ( .A(g27588), .ZN(I36454) );
INV_X32 U_g27981 ( .A(I36454), .ZN(g27981) );
INV_X32 U_I36459 ( .A(g27258), .ZN(I36459) );
INV_X32 U_g27986 ( .A(I36459), .ZN(g27986) );
INV_X32 U_I36462 ( .A(g27259), .ZN(I36462) );
INV_X32 U_g27987 ( .A(I36462), .ZN(g27987) );
INV_X32 U_I36465 ( .A(g27260), .ZN(I36465) );
INV_X32 U_g27988 ( .A(I36465), .ZN(g27988) );
INV_X32 U_I36468 ( .A(g27261), .ZN(I36468) );
INV_X32 U_g27989 ( .A(I36468), .ZN(g27989) );
INV_X32 U_g27990 ( .A(g27367), .ZN(g27990) );
INV_X32 U_I36473 ( .A(g27262), .ZN(I36473) );
INV_X32 U_g27992 ( .A(I36473), .ZN(g27992) );
INV_X32 U_I36476 ( .A(g27263), .ZN(I36476) );
INV_X32 U_g27993 ( .A(I36476), .ZN(g27993) );
INV_X32 U_I36479 ( .A(g27504), .ZN(I36479) );
INV_X32 U_g27994 ( .A(I36479), .ZN(g27994) );
INV_X32 U_I36483 ( .A(g27264), .ZN(I36483) );
INV_X32 U_g27998 ( .A(I36483), .ZN(g27998) );
INV_X32 U_I36486 ( .A(g27507), .ZN(I36486) );
INV_X32 U_g27999 ( .A(I36486), .ZN(g27999) );
INV_X32 U_I36490 ( .A(g27265), .ZN(I36490) );
INV_X32 U_g28003 ( .A(I36490), .ZN(g28003) );
INV_X32 U_I36493 ( .A(g27266), .ZN(I36493) );
INV_X32 U_g28004 ( .A(I36493), .ZN(g28004) );
INV_X32 U_I36496 ( .A(g27267), .ZN(I36496) );
INV_X32 U_g28005 ( .A(I36496), .ZN(g28005) );
INV_X32 U_I36499 ( .A(g27268), .ZN(I36499) );
INV_X32 U_g28006 ( .A(I36499), .ZN(g28006) );
INV_X32 U_I36502 ( .A(g27269), .ZN(I36502) );
INV_X32 U_g28007 ( .A(I36502), .ZN(g28007) );
INV_X32 U_I36507 ( .A(g27270), .ZN(I36507) );
INV_X32 U_g28010 ( .A(I36507), .ZN(g28010) );
INV_X32 U_I36510 ( .A(g27271), .ZN(I36510) );
INV_X32 U_g28011 ( .A(I36510), .ZN(g28011) );
INV_X32 U_I36513 ( .A(g27272), .ZN(I36513) );
INV_X32 U_g28012 ( .A(I36513), .ZN(g28012) );
INV_X32 U_I36516 ( .A(g27273), .ZN(I36516) );
INV_X32 U_g28013 ( .A(I36516), .ZN(g28013) );
INV_X32 U_g28014 ( .A(g27373), .ZN(g28014) );
INV_X32 U_I36521 ( .A(g27274), .ZN(I36521) );
INV_X32 U_g28016 ( .A(I36521), .ZN(g28016) );
INV_X32 U_I36524 ( .A(g27275), .ZN(I36524) );
INV_X32 U_g28017 ( .A(I36524), .ZN(g28017) );
INV_X32 U_I36527 ( .A(g27524), .ZN(I36527) );
INV_X32 U_g28018 ( .A(I36527), .ZN(g28018) );
INV_X32 U_I36530 ( .A(g27276), .ZN(I36530) );
INV_X32 U_g28021 ( .A(I36530), .ZN(g28021) );
INV_X32 U_I36533 ( .A(g27277), .ZN(I36533) );
INV_X32 U_g28022 ( .A(I36533), .ZN(g28022) );
INV_X32 U_I36536 ( .A(g27278), .ZN(I36536) );
INV_X32 U_g28023 ( .A(I36536), .ZN(g28023) );
INV_X32 U_I36539 ( .A(g27279), .ZN(I36539) );
INV_X32 U_g28024 ( .A(I36539), .ZN(g28024) );
INV_X32 U_I36542 ( .A(g27280), .ZN(I36542) );
INV_X32 U_g28025 ( .A(I36542), .ZN(g28025) );
INV_X32 U_I36545 ( .A(g27281), .ZN(I36545) );
INV_X32 U_g28026 ( .A(I36545), .ZN(g28026) );
INV_X32 U_I36551 ( .A(g27282), .ZN(I36551) );
INV_X32 U_g28030 ( .A(I36551), .ZN(g28030) );
INV_X32 U_I36554 ( .A(g27283), .ZN(I36554) );
INV_X32 U_g28031 ( .A(I36554), .ZN(g28031) );
INV_X32 U_I36557 ( .A(g27284), .ZN(I36557) );
INV_X32 U_g28032 ( .A(I36557), .ZN(g28032) );
INV_X32 U_I36560 ( .A(g27285), .ZN(I36560) );
INV_X32 U_g28033 ( .A(I36560), .ZN(g28033) );
INV_X32 U_I36563 ( .A(g27286), .ZN(I36563) );
INV_X32 U_g28034 ( .A(I36563), .ZN(g28034) );
INV_X32 U_I36568 ( .A(g27287), .ZN(I36568) );
INV_X32 U_g28037 ( .A(I36568), .ZN(g28037) );
INV_X32 U_I36571 ( .A(g27288), .ZN(I36571) );
INV_X32 U_g28038 ( .A(I36571), .ZN(g28038) );
INV_X32 U_I36574 ( .A(g27289), .ZN(I36574) );
INV_X32 U_g28039 ( .A(I36574), .ZN(g28039) );
INV_X32 U_I36577 ( .A(g27290), .ZN(I36577) );
INV_X32 U_g28040 ( .A(I36577), .ZN(g28040) );
INV_X32 U_g28041 ( .A(g27376), .ZN(g28041) );
INV_X32 U_I36582 ( .A(g27291), .ZN(I36582) );
INV_X32 U_g28043 ( .A(I36582), .ZN(g28043) );
INV_X32 U_I36585 ( .A(g27292), .ZN(I36585) );
INV_X32 U_g28044 ( .A(I36585), .ZN(g28044) );
INV_X32 U_I36588 ( .A(g27293), .ZN(I36588) );
INV_X32 U_g28045 ( .A(I36588), .ZN(g28045) );
INV_X32 U_I36598 ( .A(g27294), .ZN(I36598) );
INV_X32 U_g28047 ( .A(I36598), .ZN(g28047) );
INV_X32 U_I36601 ( .A(g27295), .ZN(I36601) );
INV_X32 U_g28048 ( .A(I36601), .ZN(g28048) );
INV_X32 U_I36604 ( .A(g27296), .ZN(I36604) );
INV_X32 U_g28049 ( .A(I36604), .ZN(g28049) );
INV_X32 U_I36609 ( .A(g27297), .ZN(I36609) );
INV_X32 U_g28052 ( .A(I36609), .ZN(g28052) );
INV_X32 U_I36612 ( .A(g27298), .ZN(I36612) );
INV_X32 U_g28053 ( .A(I36612), .ZN(g28053) );
INV_X32 U_I36615 ( .A(g27299), .ZN(I36615) );
INV_X32 U_g28054 ( .A(I36615), .ZN(g28054) );
INV_X32 U_I36618 ( .A(g27300), .ZN(I36618) );
INV_X32 U_g28055 ( .A(I36618), .ZN(g28055) );
INV_X32 U_I36621 ( .A(g27301), .ZN(I36621) );
INV_X32 U_g28056 ( .A(I36621), .ZN(g28056) );
INV_X32 U_I36627 ( .A(g27302), .ZN(I36627) );
INV_X32 U_g28060 ( .A(I36627), .ZN(g28060) );
INV_X32 U_I36630 ( .A(g27303), .ZN(I36630) );
INV_X32 U_g28061 ( .A(I36630), .ZN(g28061) );
INV_X32 U_I36633 ( .A(g27304), .ZN(I36633) );
INV_X32 U_g28062 ( .A(I36633), .ZN(g28062) );
INV_X32 U_I36636 ( .A(g27305), .ZN(I36636) );
INV_X32 U_g28063 ( .A(I36636), .ZN(g28063) );
INV_X32 U_I36639 ( .A(g27306), .ZN(I36639) );
INV_X32 U_g28064 ( .A(I36639), .ZN(g28064) );
INV_X32 U_I36644 ( .A(g27307), .ZN(I36644) );
INV_X32 U_g28067 ( .A(I36644), .ZN(g28067) );
INV_X32 U_I36647 ( .A(g27308), .ZN(I36647) );
INV_X32 U_g28068 ( .A(I36647), .ZN(g28068) );
INV_X32 U_I36650 ( .A(g27309), .ZN(I36650) );
INV_X32 U_g28069 ( .A(I36650), .ZN(g28069) );
INV_X32 U_I36653 ( .A(g27310), .ZN(I36653) );
INV_X32 U_g28070 ( .A(I36653), .ZN(g28070) );
INV_X32 U_I36656 ( .A(g27311), .ZN(I36656) );
INV_X32 U_g28071 ( .A(I36656), .ZN(g28071) );
INV_X32 U_I36659 ( .A(g27312), .ZN(I36659) );
INV_X32 U_g28072 ( .A(I36659), .ZN(g28072) );
INV_X32 U_I36663 ( .A(g27313), .ZN(I36663) );
INV_X32 U_g28074 ( .A(I36663), .ZN(g28074) );
INV_X32 U_I36673 ( .A(g27314), .ZN(I36673) );
INV_X32 U_g28076 ( .A(I36673), .ZN(g28076) );
INV_X32 U_I36676 ( .A(g27315), .ZN(I36676) );
INV_X32 U_g28077 ( .A(I36676), .ZN(g28077) );
INV_X32 U_I36679 ( .A(g27316), .ZN(I36679) );
INV_X32 U_g28078 ( .A(I36679), .ZN(g28078) );
INV_X32 U_I36684 ( .A(g27317), .ZN(I36684) );
INV_X32 U_g28081 ( .A(I36684), .ZN(g28081) );
INV_X32 U_I36687 ( .A(g27318), .ZN(I36687) );
INV_X32 U_g28082 ( .A(I36687), .ZN(g28082) );
INV_X32 U_I36690 ( .A(g27319), .ZN(I36690) );
INV_X32 U_g28083 ( .A(I36690), .ZN(g28083) );
INV_X32 U_I36693 ( .A(g27320), .ZN(I36693) );
INV_X32 U_g28084 ( .A(I36693), .ZN(g28084) );
INV_X32 U_I36696 ( .A(g27321), .ZN(I36696) );
INV_X32 U_g28085 ( .A(I36696), .ZN(g28085) );
INV_X32 U_I36702 ( .A(g27322), .ZN(I36702) );
INV_X32 U_g28089 ( .A(I36702), .ZN(g28089) );
INV_X32 U_I36705 ( .A(g27323), .ZN(I36705) );
INV_X32 U_g28090 ( .A(I36705), .ZN(g28090) );
INV_X32 U_I36708 ( .A(g27324), .ZN(I36708) );
INV_X32 U_g28091 ( .A(I36708), .ZN(g28091) );
INV_X32 U_I36711 ( .A(g27325), .ZN(I36711) );
INV_X32 U_g28092 ( .A(I36711), .ZN(g28092) );
INV_X32 U_I36714 ( .A(g27326), .ZN(I36714) );
INV_X32 U_g28093 ( .A(I36714), .ZN(g28093) );
INV_X32 U_I36718 ( .A(g27327), .ZN(I36718) );
INV_X32 U_g28095 ( .A(I36718), .ZN(g28095) );
INV_X32 U_I36721 ( .A(g27328), .ZN(I36721) );
INV_X32 U_g28096 ( .A(I36721), .ZN(g28096) );
INV_X32 U_I36724 ( .A(g27329), .ZN(I36724) );
INV_X32 U_g28097 ( .A(I36724), .ZN(g28097) );
INV_X32 U_I36728 ( .A(g27330), .ZN(I36728) );
INV_X32 U_g28099 ( .A(I36728), .ZN(g28099) );
INV_X32 U_I36738 ( .A(g27331), .ZN(I36738) );
INV_X32 U_g28101 ( .A(I36738), .ZN(g28101) );
INV_X32 U_I36741 ( .A(g27332), .ZN(I36741) );
INV_X32 U_g28102 ( .A(I36741), .ZN(g28102) );
INV_X32 U_I36744 ( .A(g27333), .ZN(I36744) );
INV_X32 U_g28103 ( .A(I36744), .ZN(g28103) );
INV_X32 U_I36749 ( .A(g27334), .ZN(I36749) );
INV_X32 U_g28106 ( .A(I36749), .ZN(g28106) );
INV_X32 U_I36752 ( .A(g27335), .ZN(I36752) );
INV_X32 U_g28107 ( .A(I36752), .ZN(g28107) );
INV_X32 U_I36755 ( .A(g27336), .ZN(I36755) );
INV_X32 U_g28108 ( .A(I36755), .ZN(g28108) );
INV_X32 U_I36758 ( .A(g27337), .ZN(I36758) );
INV_X32 U_g28109 ( .A(I36758), .ZN(g28109) );
INV_X32 U_I36761 ( .A(g27338), .ZN(I36761) );
INV_X32 U_g28110 ( .A(I36761), .ZN(g28110) );
INV_X32 U_I36766 ( .A(g27339), .ZN(I36766) );
INV_X32 U_g28113 ( .A(I36766), .ZN(g28113) );
INV_X32 U_I36769 ( .A(g27340), .ZN(I36769) );
INV_X32 U_g28114 ( .A(I36769), .ZN(g28114) );
INV_X32 U_I36772 ( .A(g27341), .ZN(I36772) );
INV_X32 U_g28115 ( .A(I36772), .ZN(g28115) );
INV_X32 U_I36776 ( .A(g27342), .ZN(I36776) );
INV_X32 U_g28117 ( .A(I36776), .ZN(g28117) );
INV_X32 U_I36786 ( .A(g27343), .ZN(I36786) );
INV_X32 U_g28119 ( .A(I36786), .ZN(g28119) );
INV_X32 U_I36789 ( .A(g27344), .ZN(I36789) );
INV_X32 U_g28120 ( .A(I36789), .ZN(g28120) );
INV_X32 U_I36792 ( .A(g27345), .ZN(I36792) );
INV_X32 U_g28121 ( .A(I36792), .ZN(g28121) );
INV_X32 U_I36797 ( .A(g27346), .ZN(I36797) );
INV_X32 U_g28124 ( .A(I36797), .ZN(g28124) );
INV_X32 U_I36800 ( .A(g27347), .ZN(I36800) );
INV_X32 U_g28125 ( .A(I36800), .ZN(g28125) );
INV_X32 U_I36803 ( .A(g27348), .ZN(I36803) );
INV_X32 U_g28126 ( .A(I36803), .ZN(g28126) );
INV_X32 U_g28128 ( .A(g27528), .ZN(g28128) );
INV_X32 U_I36808 ( .A(g27354), .ZN(I36808) );
INV_X32 U_g28132 ( .A(I36808), .ZN(g28132) );
INV_X32 U_g28133 ( .A(g27550), .ZN(g28133) );
INV_X32 U_g28137 ( .A(g27566), .ZN(g28137) );
INV_X32 U_g28141 ( .A(g27576), .ZN(g28141) );
INV_X32 U_g28149 ( .A(g27667), .ZN(g28149) );
INV_X32 U_g28150 ( .A(g27387), .ZN(g28150) );
INV_X32 U_g28151 ( .A(g27381), .ZN(g28151) );
INV_X32 U_g28152 ( .A(g27391), .ZN(g28152) );
INV_X32 U_g28153 ( .A(g27397), .ZN(g28153) );
INV_X32 U_g28154 ( .A(g27401), .ZN(g28154) );
INV_X32 U_g28155 ( .A(g27404), .ZN(g28155) );
INV_X32 U_g28156 ( .A(g27410), .ZN(g28156) );
INV_X32 U_g28158 ( .A(g27416), .ZN(g28158) );
INV_X32 U_g28159 ( .A(g27419), .ZN(g28159) );
INV_X32 U_g28160 ( .A(g27422), .ZN(g28160) );
INV_X32 U_g28161 ( .A(g27428), .ZN(g28161) );
INV_X32 U_g28162 ( .A(g27432), .ZN(g28162) );
INV_X32 U_g28163 ( .A(g27437), .ZN(g28163) );
INV_X32 U_g28164 ( .A(g27440), .ZN(g28164) );
INV_X32 U_g28165 ( .A(g27443), .ZN(g28165) );
INV_X32 U_g28166 ( .A(g27451), .ZN(g28166) );
INV_X32 U_g28167 ( .A(g27456), .ZN(g28167) );
INV_X32 U_g28168 ( .A(g27459), .ZN(g28168) );
INV_X32 U_g28169 ( .A(g27467), .ZN(g28169) );
INV_X32 U_g28170 ( .A(g27472), .ZN(g28170) );
INV_X32 U_g28172 ( .A(g27475), .ZN(g28172) );
INV_X32 U_g28173 ( .A(g27486), .ZN(g28173) );
INV_X32 U_g28174 ( .A(g27489), .ZN(g28174) );
INV_X32 U_g28175 ( .A(g27498), .ZN(g28175) );
INV_X32 U_g28177 ( .A(g27510), .ZN(g28177) );
INV_X32 U_g28178 ( .A(g27518), .ZN(g28178) );
INV_X32 U_I36848 ( .A(g27383), .ZN(I36848) );
INV_X32 U_g28179 ( .A(I36848), .ZN(g28179) );
INV_X32 U_g28186 ( .A(g27535), .ZN(g28186) );
INV_X32 U_g28187 ( .A(g27543), .ZN(g28187) );
INV_X32 U_g28190 ( .A(g27555), .ZN(g28190) );
INV_X32 U_I36860 ( .A(g27386), .ZN(I36860) );
INV_X32 U_g28194 ( .A(I36860), .ZN(g28194) );
INV_X32 U_I36864 ( .A(g27384), .ZN(I36864) );
INV_X32 U_g28200 ( .A(I36864), .ZN(g28200) );
INV_X32 U_I36867 ( .A(g27786), .ZN(I36867) );
INV_X32 U_g28206 ( .A(I36867), .ZN(g28206) );
INV_X32 U_I36870 ( .A(g27955), .ZN(I36870) );
INV_X32 U_g28207 ( .A(I36870), .ZN(g28207) );
INV_X32 U_I36873 ( .A(g27971), .ZN(I36873) );
INV_X32 U_g28208 ( .A(I36873), .ZN(g28208) );
INV_X32 U_I36876 ( .A(g27986), .ZN(I36876) );
INV_X32 U_g28209 ( .A(I36876), .ZN(g28209) );
INV_X32 U_I36879 ( .A(g27972), .ZN(I36879) );
INV_X32 U_g28210 ( .A(I36879), .ZN(g28210) );
INV_X32 U_I36882 ( .A(g27987), .ZN(I36882) );
INV_X32 U_g28211 ( .A(I36882), .ZN(g28211) );
INV_X32 U_I36885 ( .A(g28003), .ZN(I36885) );
INV_X32 U_g28212 ( .A(I36885), .ZN(g28212) );
INV_X32 U_I36888 ( .A(g27988), .ZN(I36888) );
INV_X32 U_g28213 ( .A(I36888), .ZN(g28213) );
INV_X32 U_I36891 ( .A(g28004), .ZN(I36891) );
INV_X32 U_g28214 ( .A(I36891), .ZN(g28214) );
INV_X32 U_I36894 ( .A(g28022), .ZN(I36894) );
INV_X32 U_g28215 ( .A(I36894), .ZN(g28215) );
INV_X32 U_I36897 ( .A(g28005), .ZN(I36897) );
INV_X32 U_g28216 ( .A(I36897), .ZN(g28216) );
INV_X32 U_I36900 ( .A(g28023), .ZN(I36900) );
INV_X32 U_g28217 ( .A(I36900), .ZN(g28217) );
INV_X32 U_I36903 ( .A(g28045), .ZN(I36903) );
INV_X32 U_g28218 ( .A(I36903), .ZN(g28218) );
INV_X32 U_I36906 ( .A(g27989), .ZN(I36906) );
INV_X32 U_g28219 ( .A(I36906), .ZN(g28219) );
INV_X32 U_I36909 ( .A(g28006), .ZN(I36909) );
INV_X32 U_g28220 ( .A(I36909), .ZN(g28220) );
INV_X32 U_I36912 ( .A(g28024), .ZN(I36912) );
INV_X32 U_g28221 ( .A(I36912), .ZN(g28221) );
INV_X32 U_I36915 ( .A(g28007), .ZN(I36915) );
INV_X32 U_g28222 ( .A(I36915), .ZN(g28222) );
INV_X32 U_I36918 ( .A(g28025), .ZN(I36918) );
INV_X32 U_g28223 ( .A(I36918), .ZN(g28223) );
INV_X32 U_I36921 ( .A(g28047), .ZN(I36921) );
INV_X32 U_g28224 ( .A(I36921), .ZN(g28224) );
INV_X32 U_I36924 ( .A(g28026), .ZN(I36924) );
INV_X32 U_g28225 ( .A(I36924), .ZN(g28225) );
INV_X32 U_I36927 ( .A(g28048), .ZN(I36927) );
INV_X32 U_g28226 ( .A(I36927), .ZN(g28226) );
INV_X32 U_I36930 ( .A(g28071), .ZN(I36930) );
INV_X32 U_g28227 ( .A(I36930), .ZN(g28227) );
INV_X32 U_I36933 ( .A(g28049), .ZN(I36933) );
INV_X32 U_g28228 ( .A(I36933), .ZN(g28228) );
INV_X32 U_I36936 ( .A(g28072), .ZN(I36936) );
INV_X32 U_g28229 ( .A(I36936), .ZN(g28229) );
INV_X32 U_I36939 ( .A(g28095), .ZN(I36939) );
INV_X32 U_g28230 ( .A(I36939), .ZN(g28230) );
INV_X32 U_I36942 ( .A(g27905), .ZN(I36942) );
INV_X32 U_g28231 ( .A(I36942), .ZN(g28231) );
INV_X32 U_I36945 ( .A(g27793), .ZN(I36945) );
INV_X32 U_g28232 ( .A(I36945), .ZN(g28232) );
INV_X32 U_I36948 ( .A(g27976), .ZN(I36948) );
INV_X32 U_g28233 ( .A(I36948), .ZN(g28233) );
INV_X32 U_I36951 ( .A(g27992), .ZN(I36951) );
INV_X32 U_g28234 ( .A(I36951), .ZN(g28234) );
INV_X32 U_I36954 ( .A(g28010), .ZN(I36954) );
INV_X32 U_g28235 ( .A(I36954), .ZN(g28235) );
INV_X32 U_I36957 ( .A(g27993), .ZN(I36957) );
INV_X32 U_g28236 ( .A(I36957), .ZN(g28236) );
INV_X32 U_I36960 ( .A(g28011), .ZN(I36960) );
INV_X32 U_g28237 ( .A(I36960), .ZN(g28237) );
INV_X32 U_I36963 ( .A(g28030), .ZN(I36963) );
INV_X32 U_g28238 ( .A(I36963), .ZN(g28238) );
INV_X32 U_I36966 ( .A(g28012), .ZN(I36966) );
INV_X32 U_g28239 ( .A(I36966), .ZN(g28239) );
INV_X32 U_I36969 ( .A(g28031), .ZN(I36969) );
INV_X32 U_g28240 ( .A(I36969), .ZN(g28240) );
INV_X32 U_I36972 ( .A(g28052), .ZN(I36972) );
INV_X32 U_g28241 ( .A(I36972), .ZN(g28241) );
INV_X32 U_I36975 ( .A(g28032), .ZN(I36975) );
INV_X32 U_g28242 ( .A(I36975), .ZN(g28242) );
INV_X32 U_I36978 ( .A(g28053), .ZN(I36978) );
INV_X32 U_g28243 ( .A(I36978), .ZN(g28243) );
INV_X32 U_I36981 ( .A(g28074), .ZN(I36981) );
INV_X32 U_g28244 ( .A(I36981), .ZN(g28244) );
INV_X32 U_I36984 ( .A(g28013), .ZN(I36984) );
INV_X32 U_g28245 ( .A(I36984), .ZN(g28245) );
INV_X32 U_I36987 ( .A(g28033), .ZN(I36987) );
INV_X32 U_g28246 ( .A(I36987), .ZN(g28246) );
INV_X32 U_I36990 ( .A(g28054), .ZN(I36990) );
INV_X32 U_g28247 ( .A(I36990), .ZN(g28247) );
INV_X32 U_I36993 ( .A(g28034), .ZN(I36993) );
INV_X32 U_g28248 ( .A(I36993), .ZN(g28248) );
INV_X32 U_I36996 ( .A(g28055), .ZN(I36996) );
INV_X32 U_g28249 ( .A(I36996), .ZN(g28249) );
INV_X32 U_I36999 ( .A(g28076), .ZN(I36999) );
INV_X32 U_g28250 ( .A(I36999), .ZN(g28250) );
INV_X32 U_I37002 ( .A(g28056), .ZN(I37002) );
INV_X32 U_g28251 ( .A(I37002), .ZN(g28251) );
INV_X32 U_I37005 ( .A(g28077), .ZN(I37005) );
INV_X32 U_g28252 ( .A(I37005), .ZN(g28252) );
INV_X32 U_I37008 ( .A(g28096), .ZN(I37008) );
INV_X32 U_g28253 ( .A(I37008), .ZN(g28253) );
INV_X32 U_I37011 ( .A(g28078), .ZN(I37011) );
INV_X32 U_g28254 ( .A(I37011), .ZN(g28254) );
INV_X32 U_I37014 ( .A(g28097), .ZN(I37014) );
INV_X32 U_g28255 ( .A(I37014), .ZN(g28255) );
INV_X32 U_I37017 ( .A(g28113), .ZN(I37017) );
INV_X32 U_g28256 ( .A(I37017), .ZN(g28256) );
INV_X32 U_I37020 ( .A(g27910), .ZN(I37020) );
INV_X32 U_g28257 ( .A(I37020), .ZN(g28257) );
INV_X32 U_I37023 ( .A(g27799), .ZN(I37023) );
INV_X32 U_g28258 ( .A(I37023), .ZN(g28258) );
INV_X32 U_I37026 ( .A(g27998), .ZN(I37026) );
INV_X32 U_g28259 ( .A(I37026), .ZN(g28259) );
INV_X32 U_I37029 ( .A(g28016), .ZN(I37029) );
INV_X32 U_g28260 ( .A(I37029), .ZN(g28260) );
INV_X32 U_I37032 ( .A(g28037), .ZN(I37032) );
INV_X32 U_g28261 ( .A(I37032), .ZN(g28261) );
INV_X32 U_I37035 ( .A(g28017), .ZN(I37035) );
INV_X32 U_g28262 ( .A(I37035), .ZN(g28262) );
INV_X32 U_I37038 ( .A(g28038), .ZN(I37038) );
INV_X32 U_g28263 ( .A(I37038), .ZN(g28263) );
INV_X32 U_I37041 ( .A(g28060), .ZN(I37041) );
INV_X32 U_g28264 ( .A(I37041), .ZN(g28264) );
INV_X32 U_I37044 ( .A(g28039), .ZN(I37044) );
INV_X32 U_g28265 ( .A(I37044), .ZN(g28265) );
INV_X32 U_I37047 ( .A(g28061), .ZN(I37047) );
INV_X32 U_g28266 ( .A(I37047), .ZN(g28266) );
INV_X32 U_I37050 ( .A(g28081), .ZN(I37050) );
INV_X32 U_g28267 ( .A(I37050), .ZN(g28267) );
INV_X32 U_I37053 ( .A(g28062), .ZN(I37053) );
INV_X32 U_g28268 ( .A(I37053), .ZN(g28268) );
INV_X32 U_I37056 ( .A(g28082), .ZN(I37056) );
INV_X32 U_g28269 ( .A(I37056), .ZN(g28269) );
INV_X32 U_I37059 ( .A(g28099), .ZN(I37059) );
INV_X32 U_g28270 ( .A(I37059), .ZN(g28270) );
INV_X32 U_I37062 ( .A(g28040), .ZN(I37062) );
INV_X32 U_g28271 ( .A(I37062), .ZN(g28271) );
INV_X32 U_I37065 ( .A(g28063), .ZN(I37065) );
INV_X32 U_g28272 ( .A(I37065), .ZN(g28272) );
INV_X32 U_I37068 ( .A(g28083), .ZN(I37068) );
INV_X32 U_g28273 ( .A(I37068), .ZN(g28273) );
INV_X32 U_I37071 ( .A(g28064), .ZN(I37071) );
INV_X32 U_g28274 ( .A(I37071), .ZN(g28274) );
INV_X32 U_I37074 ( .A(g28084), .ZN(I37074) );
INV_X32 U_g28275 ( .A(I37074), .ZN(g28275) );
INV_X32 U_I37077 ( .A(g28101), .ZN(I37077) );
INV_X32 U_g28276 ( .A(I37077), .ZN(g28276) );
INV_X32 U_I37080 ( .A(g28085), .ZN(I37080) );
INV_X32 U_g28277 ( .A(I37080), .ZN(g28277) );
INV_X32 U_I37083 ( .A(g28102), .ZN(I37083) );
INV_X32 U_g28278 ( .A(I37083), .ZN(g28278) );
INV_X32 U_I37086 ( .A(g28114), .ZN(I37086) );
INV_X32 U_g28279 ( .A(I37086), .ZN(g28279) );
INV_X32 U_I37089 ( .A(g28103), .ZN(I37089) );
INV_X32 U_g28280 ( .A(I37089), .ZN(g28280) );
INV_X32 U_I37092 ( .A(g28115), .ZN(I37092) );
INV_X32 U_g28281 ( .A(I37092), .ZN(g28281) );
INV_X32 U_I37095 ( .A(g28124), .ZN(I37095) );
INV_X32 U_g28282 ( .A(I37095), .ZN(g28282) );
INV_X32 U_I37098 ( .A(g27918), .ZN(I37098) );
INV_X32 U_g28283 ( .A(I37098), .ZN(g28283) );
INV_X32 U_I37101 ( .A(g27805), .ZN(I37101) );
INV_X32 U_g28284 ( .A(I37101), .ZN(g28284) );
INV_X32 U_I37104 ( .A(g28021), .ZN(I37104) );
INV_X32 U_g28285 ( .A(I37104), .ZN(g28285) );
INV_X32 U_I37107 ( .A(g28043), .ZN(I37107) );
INV_X32 U_g28286 ( .A(I37107), .ZN(g28286) );
INV_X32 U_I37110 ( .A(g28067), .ZN(I37110) );
INV_X32 U_g28287 ( .A(I37110), .ZN(g28287) );
INV_X32 U_I37113 ( .A(g28044), .ZN(I37113) );
INV_X32 U_g28288 ( .A(I37113), .ZN(g28288) );
INV_X32 U_I37116 ( .A(g28068), .ZN(I37116) );
INV_X32 U_g28289 ( .A(I37116), .ZN(g28289) );
INV_X32 U_I37119 ( .A(g28089), .ZN(I37119) );
INV_X32 U_g28290 ( .A(I37119), .ZN(g28290) );
INV_X32 U_I37122 ( .A(g28069), .ZN(I37122) );
INV_X32 U_g28291 ( .A(I37122), .ZN(g28291) );
INV_X32 U_I37125 ( .A(g28090), .ZN(I37125) );
INV_X32 U_g28292 ( .A(I37125), .ZN(g28292) );
INV_X32 U_I37128 ( .A(g28106), .ZN(I37128) );
INV_X32 U_g28293 ( .A(I37128), .ZN(g28293) );
INV_X32 U_I37131 ( .A(g28091), .ZN(I37131) );
INV_X32 U_g28294 ( .A(I37131), .ZN(g28294) );
INV_X32 U_I37134 ( .A(g28107), .ZN(I37134) );
INV_X32 U_g28295 ( .A(I37134), .ZN(g28295) );
INV_X32 U_I37137 ( .A(g28117), .ZN(I37137) );
INV_X32 U_g28296 ( .A(I37137), .ZN(g28296) );
INV_X32 U_I37140 ( .A(g28070), .ZN(I37140) );
INV_X32 U_g28297 ( .A(I37140), .ZN(g28297) );
INV_X32 U_I37143 ( .A(g28092), .ZN(I37143) );
INV_X32 U_g28298 ( .A(I37143), .ZN(g28298) );
INV_X32 U_I37146 ( .A(g28108), .ZN(I37146) );
INV_X32 U_g28299 ( .A(I37146), .ZN(g28299) );
INV_X32 U_I37149 ( .A(g28093), .ZN(I37149) );
INV_X32 U_g28300 ( .A(I37149), .ZN(g28300) );
INV_X32 U_I37152 ( .A(g28109), .ZN(I37152) );
INV_X32 U_g28301 ( .A(I37152), .ZN(g28301) );
INV_X32 U_I37155 ( .A(g28119), .ZN(I37155) );
INV_X32 U_g28302 ( .A(I37155), .ZN(g28302) );
INV_X32 U_I37158 ( .A(g28110), .ZN(I37158) );
INV_X32 U_g28303 ( .A(I37158), .ZN(g28303) );
INV_X32 U_I37161 ( .A(g28120), .ZN(I37161) );
INV_X32 U_g28304 ( .A(I37161), .ZN(g28304) );
INV_X32 U_I37164 ( .A(g28125), .ZN(I37164) );
INV_X32 U_g28305 ( .A(I37164), .ZN(g28305) );
INV_X32 U_I37167 ( .A(g28121), .ZN(I37167) );
INV_X32 U_g28306 ( .A(I37167), .ZN(g28306) );
INV_X32 U_I37170 ( .A(g28126), .ZN(I37170) );
INV_X32 U_g28307 ( .A(I37170), .ZN(g28307) );
INV_X32 U_I37173 ( .A(g28132), .ZN(I37173) );
INV_X32 U_g28308 ( .A(I37173), .ZN(g28308) );
INV_X32 U_I37176 ( .A(g27927), .ZN(I37176) );
INV_X32 U_g28309 ( .A(I37176), .ZN(g28309) );
INV_X32 U_I37179 ( .A(g27784), .ZN(I37179) );
INV_X32 U_g28310 ( .A(I37179), .ZN(g28310) );
INV_X32 U_I37182 ( .A(g27791), .ZN(I37182) );
INV_X32 U_g28311 ( .A(I37182), .ZN(g28311) );
INV_X32 U_I37185 ( .A(g27797), .ZN(I37185) );
INV_X32 U_g28312 ( .A(I37185), .ZN(g28312) );
INV_X32 U_I37188 ( .A(g27785), .ZN(I37188) );
INV_X32 U_g28313 ( .A(I37188), .ZN(g28313) );
INV_X32 U_I37191 ( .A(g27792), .ZN(I37191) );
INV_X32 U_g28314 ( .A(I37191), .ZN(g28314) );
INV_X32 U_I37194 ( .A(g27800), .ZN(I37194) );
INV_X32 U_g28315 ( .A(I37194), .ZN(g28315) );
INV_X32 U_I37197 ( .A(g27903), .ZN(I37197) );
INV_X32 U_g28316 ( .A(I37197), .ZN(g28316) );
INV_X32 U_I37200 ( .A(g27907), .ZN(I37200) );
INV_X32 U_g28317 ( .A(I37200), .ZN(g28317) );
INV_X32 U_I37203 ( .A(g27912), .ZN(I37203) );
INV_X32 U_g28318 ( .A(I37203), .ZN(g28318) );
INV_X32 U_I37228 ( .A(g28194), .ZN(I37228) );
INV_X32 U_g28341 ( .A(I37228), .ZN(g28341) );
INV_X32 U_I37232 ( .A(g28200), .ZN(I37232) );
INV_X32 U_g28343 ( .A(I37232), .ZN(g28343) );
INV_X32 U_I37238 ( .A(g28179), .ZN(I37238) );
INV_X32 U_g28347 ( .A(I37238), .ZN(g28347) );
INV_X32 U_I37252 ( .A(g28200), .ZN(I37252) );
INV_X32 U_g28359 ( .A(I37252), .ZN(g28359) );
INV_X32 U_I37260 ( .A(g28179), .ZN(I37260) );
INV_X32 U_g28365 ( .A(I37260), .ZN(g28365) );
INV_X32 U_I37266 ( .A(g28200), .ZN(I37266) );
INV_X32 U_g28369 ( .A(I37266), .ZN(g28369) );
INV_X32 U_I37269 ( .A(g28145), .ZN(I37269) );
INV_X32 U_g28370 ( .A(I37269), .ZN(g28370) );
INV_X32 U_I37273 ( .A(g28179), .ZN(I37273) );
INV_X32 U_g28372 ( .A(I37273), .ZN(g28372) );
INV_X32 U_I37277 ( .A(g28146), .ZN(I37277) );
INV_X32 U_g28374 ( .A(I37277), .ZN(g28374) );
INV_X32 U_I37280 ( .A(g28179), .ZN(I37280) );
INV_X32 U_g28375 ( .A(I37280), .ZN(g28375) );
INV_X32 U_I37284 ( .A(g28147), .ZN(I37284) );
INV_X32 U_g28377 ( .A(I37284), .ZN(g28377) );
INV_X32 U_I37291 ( .A(g28148), .ZN(I37291) );
INV_X32 U_g28382 ( .A(I37291), .ZN(g28382) );
INV_X32 U_I37319 ( .A(g28149), .ZN(I37319) );
INV_X32 U_g28390 ( .A(I37319), .ZN(g28390) );
INV_X32 U_I37330 ( .A(g28194), .ZN(I37330) );
INV_X32 U_g28393 ( .A(I37330), .ZN(g28393) );
INV_X32 U_I37334 ( .A(g28194), .ZN(I37334) );
INV_X32 U_g28395 ( .A(I37334), .ZN(g28395) );
INV_X32 U_g28419 ( .A(g28151), .ZN(g28419) );
INV_X32 U_I37379 ( .A(g28199), .ZN(I37379) );
INV_X32 U_g28432 ( .A(I37379), .ZN(g28432) );
INV_X32 U_I37386 ( .A(g28194), .ZN(I37386) );
INV_X32 U_g28437 ( .A(I37386), .ZN(g28437) );
INV_X32 U_I37394 ( .A(g27718), .ZN(I37394) );
INV_X32 U_g28443 ( .A(I37394), .ZN(g28443) );
INV_X32 U_I37400 ( .A(g28200), .ZN(I37400) );
INV_X32 U_g28447 ( .A(I37400), .ZN(g28447) );
INV_X32 U_I37410 ( .A(g27722), .ZN(I37410) );
INV_X32 U_g28455 ( .A(I37410), .ZN(g28455) );
INV_X32 U_I37415 ( .A(g28179), .ZN(I37415) );
INV_X32 U_g28458 ( .A(I37415), .ZN(g28458) );
INV_X32 U_I37426 ( .A(g27724), .ZN(I37426) );
INV_X32 U_g28467 ( .A(I37426), .ZN(g28467) );
INV_X32 U_g28483 ( .A(g27776), .ZN(g28483) );
INV_X32 U_g28491 ( .A(g27780), .ZN(g28491) );
INV_X32 U_g28496 ( .A(g27787), .ZN(g28496) );
INV_X32 U_I37459 ( .A(g27759), .ZN(I37459) );
INV_X32 U_g28498 ( .A(I37459), .ZN(g28498) );
INV_X32 U_g28500 ( .A(g27794), .ZN(g28500) );
INV_X32 U_I37467 ( .A(g27760), .ZN(I37467) );
INV_X32 U_g28524 ( .A(I37467), .ZN(g28524) );
INV_X32 U_I37471 ( .A(g27761), .ZN(I37471) );
INV_X32 U_g28526 ( .A(I37471), .ZN(g28526) );
INV_X32 U_I37474 ( .A(g27762), .ZN(I37474) );
INV_X32 U_g28527 ( .A(I37474), .ZN(g28527) );
INV_X32 U_I37481 ( .A(g27763), .ZN(I37481) );
INV_X32 U_g28552 ( .A(I37481), .ZN(g28552) );
INV_X32 U_I37484 ( .A(g27764), .ZN(I37484) );
INV_X32 U_g28553 ( .A(I37484), .ZN(g28553) );
INV_X32 U_g28554 ( .A(g27806), .ZN(g28554) );
INV_X32 U_I37488 ( .A(g27765), .ZN(I37488) );
INV_X32 U_g28555 ( .A(I37488), .ZN(g28555) );
INV_X32 U_I37494 ( .A(g27766), .ZN(I37494) );
INV_X32 U_g28579 ( .A(I37494), .ZN(g28579) );
INV_X32 U_I37497 ( .A(g27767), .ZN(I37497) );
INV_X32 U_g28580 ( .A(I37497), .ZN(g28580) );
INV_X32 U_g28581 ( .A(g27817), .ZN(g28581) );
INV_X32 U_g28582 ( .A(g27820), .ZN(g28582) );
INV_X32 U_I37502 ( .A(g27768), .ZN(I37502) );
INV_X32 U_g28583 ( .A(I37502), .ZN(g28583) );
INV_X32 U_I37508 ( .A(g27769), .ZN(I37508) );
INV_X32 U_g28607 ( .A(I37508), .ZN(g28607) );
INV_X32 U_g28608 ( .A(g27831), .ZN(g28608) );
INV_X32 U_g28609 ( .A(g27839), .ZN(g28609) );
INV_X32 U_g28610 ( .A(g27843), .ZN(g28610) );
INV_X32 U_I37514 ( .A(g27771), .ZN(I37514) );
INV_X32 U_g28611 ( .A(I37514), .ZN(g28611) );
INV_X32 U_g28612 ( .A(g28046), .ZN(g28612) );
INV_X32 U_g28616 ( .A(g27847), .ZN(g28616) );
INV_X32 U_g28617 ( .A(g27858), .ZN(g28617) );
INV_X32 U_g28618 ( .A(g27861), .ZN(g28618) );
INV_X32 U_g28619 ( .A(g28075), .ZN(g28619) );
INV_X32 U_g28623 ( .A(g27872), .ZN(g28623) );
INV_X32 U_g28624 ( .A(g27879), .ZN(g28624) );
INV_X32 U_g28625 ( .A(g28100), .ZN(g28625) );
INV_X32 U_g28629 ( .A(g27889), .ZN(g28629) );
INV_X32 U_g28630 ( .A(g28118), .ZN(g28630) );
INV_X32 U_g28638 ( .A(g28200), .ZN(g28638) );
INV_X32 U_g28639 ( .A(g27919), .ZN(g28639) );
INV_X32 U_g28640 ( .A(g27928), .ZN(g28640) );
INV_X32 U_g28641 ( .A(g27932), .ZN(g28641) );
INV_X32 U_g28642 ( .A(g27939), .ZN(g28642) );
INV_X32 U_g28643 ( .A(g27942), .ZN(g28643) );
INV_X32 U_g28644 ( .A(g27946), .ZN(g28644) );
INV_X32 U_g28645 ( .A(g27952), .ZN(g28645) );
INV_X32 U_g28646 ( .A(g27956), .ZN(g28646) );
INV_X32 U_g28647 ( .A(g27959), .ZN(g28647) );
INV_X32 U_g28648 ( .A(g27965), .ZN(g28648) );
INV_X32 U_g28649 ( .A(g27973), .ZN(g28649) );
INV_X32 U_g28650 ( .A(g27977), .ZN(g28650) );
INV_X32 U_g28651 ( .A(g27981), .ZN(g28651) );
INV_X32 U_g28652 ( .A(g27994), .ZN(g28652) );
INV_X32 U_g28653 ( .A(g27999), .ZN(g28653) );
INV_X32 U_g28655 ( .A(g28018), .ZN(g28655) );
INV_X32 U_I37566 ( .A(g28370), .ZN(I37566) );
INV_X32 U_g28673 ( .A(I37566), .ZN(g28673) );
INV_X32 U_I37569 ( .A(g28498), .ZN(I37569) );
INV_X32 U_g28674 ( .A(I37569), .ZN(g28674) );
INV_X32 U_I37572 ( .A(g28524), .ZN(I37572) );
INV_X32 U_g28675 ( .A(I37572), .ZN(g28675) );
INV_X32 U_I37575 ( .A(g28527), .ZN(I37575) );
INV_X32 U_g28676 ( .A(I37575), .ZN(g28676) );
INV_X32 U_I37578 ( .A(g28432), .ZN(I37578) );
INV_X32 U_g28677 ( .A(I37578), .ZN(g28677) );
INV_X32 U_I37581 ( .A(g28374), .ZN(I37581) );
INV_X32 U_g28678 ( .A(I37581), .ZN(g28678) );
INV_X32 U_I37584 ( .A(g28526), .ZN(I37584) );
INV_X32 U_g28679 ( .A(I37584), .ZN(g28679) );
INV_X32 U_I37587 ( .A(g28552), .ZN(I37587) );
INV_X32 U_g28680 ( .A(I37587), .ZN(g28680) );
INV_X32 U_I37590 ( .A(g28555), .ZN(I37590) );
INV_X32 U_g28681 ( .A(I37590), .ZN(g28681) );
INV_X32 U_I37593 ( .A(g28443), .ZN(I37593) );
INV_X32 U_g28682 ( .A(I37593), .ZN(g28682) );
INV_X32 U_I37596 ( .A(g28377), .ZN(I37596) );
INV_X32 U_g28683 ( .A(I37596), .ZN(g28683) );
INV_X32 U_I37599 ( .A(g28553), .ZN(I37599) );
INV_X32 U_g28684 ( .A(I37599), .ZN(g28684) );
INV_X32 U_I37602 ( .A(g28579), .ZN(I37602) );
INV_X32 U_g28685 ( .A(I37602), .ZN(g28685) );
INV_X32 U_I37605 ( .A(g28583), .ZN(I37605) );
INV_X32 U_g28686 ( .A(I37605), .ZN(g28686) );
INV_X32 U_I37608 ( .A(g28455), .ZN(I37608) );
INV_X32 U_g28687 ( .A(I37608), .ZN(g28687) );
INV_X32 U_I37611 ( .A(g28382), .ZN(I37611) );
INV_X32 U_g28688 ( .A(I37611), .ZN(g28688) );
INV_X32 U_I37614 ( .A(g28580), .ZN(I37614) );
INV_X32 U_g28689 ( .A(I37614), .ZN(g28689) );
INV_X32 U_I37617 ( .A(g28607), .ZN(I37617) );
INV_X32 U_g28690 ( .A(I37617), .ZN(g28690) );
INV_X32 U_I37620 ( .A(g28611), .ZN(I37620) );
INV_X32 U_g28691 ( .A(I37620), .ZN(g28691) );
INV_X32 U_I37623 ( .A(g28467), .ZN(I37623) );
INV_X32 U_g28692 ( .A(I37623), .ZN(g28692) );
INV_X32 U_I37626 ( .A(g28393), .ZN(I37626) );
INV_X32 U_g28693 ( .A(I37626), .ZN(g28693) );
INV_X32 U_I37629 ( .A(g28369), .ZN(I37629) );
INV_X32 U_g28694 ( .A(I37629), .ZN(g28694) );
INV_X32 U_I37632 ( .A(g28372), .ZN(I37632) );
INV_X32 U_g28695 ( .A(I37632), .ZN(g28695) );
INV_X32 U_I37635 ( .A(g28390), .ZN(I37635) );
INV_X32 U_g28696 ( .A(I37635), .ZN(g28696) );
INV_X32 U_I37638 ( .A(g28395), .ZN(I37638) );
INV_X32 U_g28697 ( .A(I37638), .ZN(g28697) );
INV_X32 U_I37641 ( .A(g28375), .ZN(I37641) );
INV_X32 U_g28698 ( .A(I37641), .ZN(g28698) );
INV_X32 U_I37644 ( .A(g28341), .ZN(I37644) );
INV_X32 U_g28699 ( .A(I37644), .ZN(g28699) );
INV_X32 U_I37647 ( .A(g28343), .ZN(I37647) );
INV_X32 U_g28700 ( .A(I37647), .ZN(g28700) );
INV_X32 U_I37650 ( .A(g28347), .ZN(I37650) );
INV_X32 U_g28701 ( .A(I37650), .ZN(g28701) );
INV_X32 U_I37653 ( .A(g28359), .ZN(I37653) );
INV_X32 U_g28702 ( .A(I37653), .ZN(g28702) );
INV_X32 U_I37656 ( .A(g28365), .ZN(I37656) );
INV_X32 U_g28703 ( .A(I37656), .ZN(g28703) );
INV_X32 U_I37659 ( .A(g28437), .ZN(I37659) );
INV_X32 U_g28704 ( .A(I37659), .ZN(g28704) );
INV_X32 U_I37662 ( .A(g28447), .ZN(I37662) );
INV_X32 U_g28705 ( .A(I37662), .ZN(g28705) );
INV_X32 U_I37665 ( .A(g28458), .ZN(I37665) );
INV_X32 U_g28706 ( .A(I37665), .ZN(g28706) );
INV_X32 U_g28720 ( .A(g28495), .ZN(g28720) );
INV_X32 U_g28721 ( .A(g28490), .ZN(g28721) );
INV_X32 U_g28723 ( .A(g28528), .ZN(g28723) );
INV_X32 U_g28725 ( .A(g28499), .ZN(g28725) );
INV_X32 U_g28727 ( .A(g28489), .ZN(g28727) );
INV_X32 U_g28730 ( .A(g28470), .ZN(g28730) );
INV_X32 U_g28734 ( .A(g28525), .ZN(g28734) );
INV_X32 U_g28740 ( .A(g28488), .ZN(g28740) );
INV_X32 U_I37702 ( .A(g28512), .ZN(I37702) );
INV_X32 U_g28741 ( .A(I37702), .ZN(g28741) );
INV_X32 U_I37712 ( .A(g28512), .ZN(I37712) );
INV_X32 U_g28751 ( .A(I37712), .ZN(g28751) );
INV_X32 U_I37716 ( .A(g28540), .ZN(I37716) );
INV_X32 U_g28755 ( .A(I37716), .ZN(g28755) );
INV_X32 U_I37725 ( .A(g28540), .ZN(I37725) );
INV_X32 U_g28764 ( .A(I37725), .ZN(g28764) );
INV_X32 U_I37729 ( .A(g28567), .ZN(I37729) );
INV_X32 U_g28768 ( .A(I37729), .ZN(g28768) );
INV_X32 U_I37736 ( .A(g28567), .ZN(I37736) );
INV_X32 U_g28775 ( .A(I37736), .ZN(g28775) );
INV_X32 U_I37740 ( .A(g28595), .ZN(I37740) );
INV_X32 U_g28779 ( .A(I37740), .ZN(g28779) );
INV_X32 U_I37746 ( .A(g28595), .ZN(I37746) );
INV_X32 U_g28785 ( .A(I37746), .ZN(g28785) );
INV_X32 U_I37752 ( .A(g28512), .ZN(I37752) );
INV_X32 U_g28791 ( .A(I37752), .ZN(g28791) );
INV_X32 U_I37757 ( .A(g28512), .ZN(I37757) );
INV_X32 U_g28796 ( .A(I37757), .ZN(g28796) );
INV_X32 U_I37760 ( .A(g28540), .ZN(I37760) );
INV_X32 U_g28799 ( .A(I37760), .ZN(g28799) );
INV_X32 U_I37765 ( .A(g28512), .ZN(I37765) );
INV_X32 U_g28804 ( .A(I37765), .ZN(g28804) );
INV_X32 U_I37768 ( .A(g28540), .ZN(I37768) );
INV_X32 U_g28807 ( .A(I37768), .ZN(g28807) );
INV_X32 U_I37771 ( .A(g28567), .ZN(I37771) );
INV_X32 U_g28810 ( .A(I37771), .ZN(g28810) );
INV_X32 U_I37775 ( .A(g28540), .ZN(I37775) );
INV_X32 U_g28814 ( .A(I37775), .ZN(g28814) );
INV_X32 U_I37778 ( .A(g28567), .ZN(I37778) );
INV_X32 U_g28817 ( .A(I37778), .ZN(g28817) );
INV_X32 U_I37781 ( .A(g28595), .ZN(I37781) );
INV_X32 U_g28820 ( .A(I37781), .ZN(g28820) );
INV_X32 U_I37784 ( .A(g28567), .ZN(I37784) );
INV_X32 U_g28823 ( .A(I37784), .ZN(g28823) );
INV_X32 U_I37787 ( .A(g28595), .ZN(I37787) );
INV_X32 U_g28826 ( .A(I37787), .ZN(g28826) );
INV_X32 U_I37790 ( .A(g28595), .ZN(I37790) );
INV_X32 U_g28829 ( .A(I37790), .ZN(g28829) );
INV_X32 U_I37793 ( .A(g28638), .ZN(I37793) );
INV_X32 U_g28832 ( .A(I37793), .ZN(g28832) );
INV_X32 U_I37796 ( .A(g28634), .ZN(I37796) );
INV_X32 U_g28833 ( .A(I37796), .ZN(g28833) );
INV_X32 U_I37800 ( .A(g28635), .ZN(I37800) );
INV_X32 U_g28835 ( .A(I37800), .ZN(g28835) );
INV_X32 U_I37804 ( .A(g28636), .ZN(I37804) );
INV_X32 U_g28837 ( .A(I37804), .ZN(g28837) );
INV_X32 U_I37808 ( .A(g28637), .ZN(I37808) );
INV_X32 U_g28839 ( .A(I37808), .ZN(g28839) );
INV_X32 U_g28855 ( .A(g28409), .ZN(g28855) );
INV_X32 U_g28859 ( .A(g28413), .ZN(g28859) );
INV_X32 U_g28863 ( .A(g28417), .ZN(g28863) );
INV_X32 U_g28867 ( .A(g28418), .ZN(g28867) );
INV_X32 U_I37842 ( .A(g28501), .ZN(I37842) );
INV_X32 U_g28871 ( .A(I37842), .ZN(g28871) );
INV_X32 U_I37846 ( .A(g28501), .ZN(I37846) );
INV_X32 U_g28877 ( .A(I37846), .ZN(g28877) );
INV_X32 U_I37851 ( .A(g28668), .ZN(I37851) );
INV_X32 U_g28882 ( .A(I37851), .ZN(g28882) );
INV_X32 U_I37854 ( .A(g28529), .ZN(I37854) );
INV_X32 U_g28883 ( .A(I37854), .ZN(g28883) );
INV_X32 U_I37858 ( .A(g28501), .ZN(I37858) );
INV_X32 U_g28889 ( .A(I37858), .ZN(g28889) );
INV_X32 U_I37863 ( .A(g28529), .ZN(I37863) );
INV_X32 U_g28894 ( .A(I37863), .ZN(g28894) );
INV_X32 U_I37868 ( .A(g28321), .ZN(I37868) );
INV_X32 U_g28899 ( .A(I37868), .ZN(g28899) );
INV_X32 U_I37871 ( .A(g28556), .ZN(I37871) );
INV_X32 U_g28900 ( .A(I37871), .ZN(g28900) );
INV_X32 U_I37875 ( .A(g28501), .ZN(I37875) );
INV_X32 U_g28906 ( .A(I37875), .ZN(g28906) );
INV_X32 U_I37880 ( .A(g28529), .ZN(I37880) );
INV_X32 U_g28911 ( .A(I37880), .ZN(g28911) );
INV_X32 U_I37885 ( .A(g28556), .ZN(I37885) );
INV_X32 U_g28916 ( .A(I37885), .ZN(g28916) );
INV_X32 U_I37891 ( .A(g28325), .ZN(I37891) );
INV_X32 U_g28924 ( .A(I37891), .ZN(g28924) );
INV_X32 U_I37894 ( .A(g28584), .ZN(I37894) );
INV_X32 U_g28925 ( .A(I37894), .ZN(g28925) );
INV_X32 U_I37897 ( .A(g28501), .ZN(I37897) );
INV_X32 U_g28928 ( .A(I37897), .ZN(g28928) );
INV_X32 U_I37901 ( .A(g28529), .ZN(I37901) );
INV_X32 U_g28932 ( .A(I37901), .ZN(g28932) );
INV_X32 U_I37906 ( .A(g28556), .ZN(I37906) );
INV_X32 U_g28937 ( .A(I37906), .ZN(g28937) );
INV_X32 U_I37912 ( .A(g28584), .ZN(I37912) );
INV_X32 U_g28945 ( .A(I37912), .ZN(g28945) );
INV_X32 U_I37917 ( .A(g28328), .ZN(I37917) );
INV_X32 U_g28950 ( .A(I37917), .ZN(g28950) );
INV_X32 U_I37920 ( .A(g28501), .ZN(I37920) );
INV_X32 U_g28951 ( .A(I37920), .ZN(g28951) );
INV_X32 U_I37924 ( .A(g28529), .ZN(I37924) );
INV_X32 U_g28955 ( .A(I37924), .ZN(g28955) );
INV_X32 U_I37928 ( .A(g28556), .ZN(I37928) );
INV_X32 U_g28959 ( .A(I37928), .ZN(g28959) );
INV_X32 U_I37934 ( .A(g28584), .ZN(I37934) );
INV_X32 U_g28967 ( .A(I37934), .ZN(g28967) );
INV_X32 U_I37939 ( .A(g28501), .ZN(I37939) );
INV_X32 U_g28972 ( .A(I37939), .ZN(g28972) );
INV_X32 U_I37942 ( .A(g28501), .ZN(I37942) );
INV_X32 U_g28975 ( .A(I37942), .ZN(g28975) );
INV_X32 U_I37946 ( .A(g28529), .ZN(I37946) );
INV_X32 U_g28979 ( .A(I37946), .ZN(g28979) );
INV_X32 U_I37950 ( .A(g28556), .ZN(I37950) );
INV_X32 U_g28983 ( .A(I37950), .ZN(g28983) );
INV_X32 U_I37956 ( .A(g28584), .ZN(I37956) );
INV_X32 U_g28993 ( .A(I37956), .ZN(g28993) );
INV_X32 U_I37961 ( .A(g28501), .ZN(I37961) );
INV_X32 U_g28998 ( .A(I37961), .ZN(g28998) );
INV_X32 U_I37965 ( .A(g28529), .ZN(I37965) );
INV_X32 U_g29002 ( .A(I37965), .ZN(g29002) );
INV_X32 U_I37968 ( .A(g28529), .ZN(I37968) );
INV_X32 U_g29005 ( .A(I37968), .ZN(g29005) );
INV_X32 U_I37973 ( .A(g28556), .ZN(I37973) );
INV_X32 U_g29010 ( .A(I37973), .ZN(g29010) );
INV_X32 U_I37978 ( .A(g28584), .ZN(I37978) );
INV_X32 U_g29019 ( .A(I37978), .ZN(g29019) );
INV_X32 U_I37982 ( .A(g28501), .ZN(I37982) );
INV_X32 U_g29023 ( .A(I37982), .ZN(g29023) );
INV_X32 U_I37986 ( .A(g28529), .ZN(I37986) );
INV_X32 U_g29027 ( .A(I37986), .ZN(g29027) );
INV_X32 U_I37991 ( .A(g28556), .ZN(I37991) );
INV_X32 U_g29032 ( .A(I37991), .ZN(g29032) );
INV_X32 U_I37994 ( .A(g28556), .ZN(I37994) );
INV_X32 U_g29035 ( .A(I37994), .ZN(g29035) );
INV_X32 U_I37999 ( .A(g28584), .ZN(I37999) );
INV_X32 U_g29042 ( .A(I37999), .ZN(g29042) );
INV_X32 U_I38003 ( .A(g28529), .ZN(I38003) );
INV_X32 U_g29046 ( .A(I38003), .ZN(g29046) );
INV_X32 U_I38007 ( .A(g28556), .ZN(I38007) );
INV_X32 U_g29050 ( .A(I38007), .ZN(g29050) );
INV_X32 U_I38011 ( .A(g28584), .ZN(I38011) );
INV_X32 U_g29054 ( .A(I38011), .ZN(g29054) );
INV_X32 U_I38014 ( .A(g28584), .ZN(I38014) );
INV_X32 U_g29057 ( .A(I38014), .ZN(g29057) );
INV_X32 U_I38018 ( .A(g28342), .ZN(I38018) );
INV_X32 U_g29061 ( .A(I38018), .ZN(g29061) );
INV_X32 U_I38024 ( .A(g28556), .ZN(I38024) );
INV_X32 U_g29065 ( .A(I38024), .ZN(g29065) );
INV_X32 U_I38028 ( .A(g28584), .ZN(I38028) );
INV_X32 U_g29069 ( .A(I38028), .ZN(g29069) );
INV_X32 U_I38032 ( .A(g28344), .ZN(I38032) );
INV_X32 U_g29073 ( .A(I38032), .ZN(g29073) );
INV_X32 U_I38035 ( .A(g28345), .ZN(I38035) );
INV_X32 U_g29074 ( .A(I38035), .ZN(g29074) );
INV_X32 U_I38038 ( .A(g28346), .ZN(I38038) );
INV_X32 U_g29075 ( .A(I38038), .ZN(g29075) );
INV_X32 U_I38042 ( .A(g28584), .ZN(I38042) );
INV_X32 U_g29077 ( .A(I38042), .ZN(g29077) );
INV_X32 U_I38046 ( .A(g28348), .ZN(I38046) );
INV_X32 U_g29081 ( .A(I38046), .ZN(g29081) );
INV_X32 U_I38049 ( .A(g28349), .ZN(I38049) );
INV_X32 U_g29082 ( .A(I38049), .ZN(g29082) );
INV_X32 U_I38053 ( .A(g28350), .ZN(I38053) );
INV_X32 U_g29084 ( .A(I38053), .ZN(g29084) );
INV_X32 U_I38056 ( .A(g28351), .ZN(I38056) );
INV_X32 U_g29085 ( .A(I38056), .ZN(g29085) );
INV_X32 U_I38059 ( .A(g28352), .ZN(I38059) );
INV_X32 U_g29086 ( .A(I38059), .ZN(g29086) );
INV_X32 U_I38064 ( .A(g28353), .ZN(I38064) );
INV_X32 U_g29089 ( .A(I38064), .ZN(g29089) );
INV_X32 U_I38068 ( .A(g28354), .ZN(I38068) );
INV_X32 U_g29091 ( .A(I38068), .ZN(g29091) );
INV_X32 U_I38071 ( .A(g28355), .ZN(I38071) );
INV_X32 U_g29092 ( .A(I38071), .ZN(g29092) );
INV_X32 U_I38074 ( .A(g28356), .ZN(I38074) );
INV_X32 U_g29093 ( .A(I38074), .ZN(g29093) );
INV_X32 U_I38077 ( .A(g28357), .ZN(I38077) );
INV_X32 U_g29094 ( .A(I38077), .ZN(g29094) );
INV_X32 U_I38080 ( .A(g28358), .ZN(I38080) );
INV_X32 U_g29095 ( .A(I38080), .ZN(g29095) );
INV_X32 U_I38085 ( .A(g28360), .ZN(I38085) );
INV_X32 U_g29098 ( .A(I38085), .ZN(g29098) );
INV_X32 U_I38088 ( .A(g28361), .ZN(I38088) );
INV_X32 U_g29099 ( .A(I38088), .ZN(g29099) );
INV_X32 U_I38091 ( .A(g28362), .ZN(I38091) );
INV_X32 U_g29100 ( .A(I38091), .ZN(g29100) );
INV_X32 U_I38094 ( .A(g28363), .ZN(I38094) );
INV_X32 U_g29101 ( .A(I38094), .ZN(g29101) );
INV_X32 U_I38097 ( .A(g28364), .ZN(I38097) );
INV_X32 U_g29102 ( .A(I38097), .ZN(g29102) );
INV_X32 U_I38101 ( .A(g28366), .ZN(I38101) );
INV_X32 U_g29104 ( .A(I38101), .ZN(g29104) );
INV_X32 U_I38104 ( .A(g28367), .ZN(I38104) );
INV_X32 U_g29105 ( .A(I38104), .ZN(g29105) );
INV_X32 U_I38107 ( .A(g28368), .ZN(I38107) );
INV_X32 U_g29106 ( .A(I38107), .ZN(g29106) );
INV_X32 U_I38111 ( .A(g28371), .ZN(I38111) );
INV_X32 U_g29108 ( .A(I38111), .ZN(g29108) );
INV_X32 U_I38119 ( .A(g28420), .ZN(I38119) );
INV_X32 U_g29117 ( .A(I38119), .ZN(g29117) );
INV_X32 U_I38122 ( .A(g28421), .ZN(I38122) );
INV_X32 U_g29118 ( .A(I38122), .ZN(g29118) );
INV_X32 U_I38125 ( .A(g28425), .ZN(I38125) );
INV_X32 U_g29119 ( .A(I38125), .ZN(g29119) );
INV_X32 U_I38128 ( .A(g28419), .ZN(I38128) );
INV_X32 U_g29120 ( .A(I38128), .ZN(g29120) );
INV_X32 U_I38136 ( .A(g28833), .ZN(I38136) );
INV_X32 U_g29131 ( .A(I38136), .ZN(g29131) );
INV_X32 U_I38139 ( .A(g29061), .ZN(I38139) );
INV_X32 U_g29132 ( .A(I38139), .ZN(g29132) );
INV_X32 U_I38142 ( .A(g29073), .ZN(I38142) );
INV_X32 U_g29133 ( .A(I38142), .ZN(g29133) );
INV_X32 U_I38145 ( .A(g29081), .ZN(I38145) );
INV_X32 U_g29134 ( .A(I38145), .ZN(g29134) );
INV_X32 U_I38148 ( .A(g29074), .ZN(I38148) );
INV_X32 U_g29135 ( .A(I38148), .ZN(g29135) );
INV_X32 U_I38151 ( .A(g29082), .ZN(I38151) );
INV_X32 U_g29136 ( .A(I38151), .ZN(g29136) );
INV_X32 U_I38154 ( .A(g29089), .ZN(I38154) );
INV_X32 U_g29137 ( .A(I38154), .ZN(g29137) );
INV_X32 U_I38157 ( .A(g28882), .ZN(I38157) );
INV_X32 U_g29138 ( .A(I38157), .ZN(g29138) );
INV_X32 U_I38160 ( .A(g28835), .ZN(I38160) );
INV_X32 U_g29139 ( .A(I38160), .ZN(g29139) );
INV_X32 U_I38163 ( .A(g29075), .ZN(I38163) );
INV_X32 U_g29140 ( .A(I38163), .ZN(g29140) );
INV_X32 U_I38166 ( .A(g29084), .ZN(I38166) );
INV_X32 U_g29141 ( .A(I38166), .ZN(g29141) );
INV_X32 U_I38169 ( .A(g29091), .ZN(I38169) );
INV_X32 U_g29142 ( .A(I38169), .ZN(g29142) );
INV_X32 U_I38172 ( .A(g29085), .ZN(I38172) );
INV_X32 U_g29143 ( .A(I38172), .ZN(g29143) );
INV_X32 U_I38175 ( .A(g29092), .ZN(I38175) );
INV_X32 U_g29144 ( .A(I38175), .ZN(g29144) );
INV_X32 U_I38178 ( .A(g29098), .ZN(I38178) );
INV_X32 U_g29145 ( .A(I38178), .ZN(g29145) );
INV_X32 U_I38181 ( .A(g28899), .ZN(I38181) );
INV_X32 U_g29146 ( .A(I38181), .ZN(g29146) );
INV_X32 U_I38184 ( .A(g28837), .ZN(I38184) );
INV_X32 U_g29147 ( .A(I38184), .ZN(g29147) );
INV_X32 U_I38187 ( .A(g29086), .ZN(I38187) );
INV_X32 U_g29148 ( .A(I38187), .ZN(g29148) );
INV_X32 U_I38190 ( .A(g29093), .ZN(I38190) );
INV_X32 U_g29149 ( .A(I38190), .ZN(g29149) );
INV_X32 U_I38193 ( .A(g29099), .ZN(I38193) );
INV_X32 U_g29150 ( .A(I38193), .ZN(g29150) );
INV_X32 U_I38196 ( .A(g29094), .ZN(I38196) );
INV_X32 U_g29151 ( .A(I38196), .ZN(g29151) );
INV_X32 U_I38199 ( .A(g29100), .ZN(I38199) );
INV_X32 U_g29152 ( .A(I38199), .ZN(g29152) );
INV_X32 U_I38202 ( .A(g29104), .ZN(I38202) );
INV_X32 U_g29153 ( .A(I38202), .ZN(g29153) );
INV_X32 U_I38205 ( .A(g28924), .ZN(I38205) );
INV_X32 U_g29154 ( .A(I38205), .ZN(g29154) );
INV_X32 U_I38208 ( .A(g28839), .ZN(I38208) );
INV_X32 U_g29155 ( .A(I38208), .ZN(g29155) );
INV_X32 U_I38211 ( .A(g29095), .ZN(I38211) );
INV_X32 U_g29156 ( .A(I38211), .ZN(g29156) );
INV_X32 U_I38214 ( .A(g29101), .ZN(I38214) );
INV_X32 U_g29157 ( .A(I38214), .ZN(g29157) );
INV_X32 U_I38217 ( .A(g29105), .ZN(I38217) );
INV_X32 U_g29158 ( .A(I38217), .ZN(g29158) );
INV_X32 U_I38220 ( .A(g29102), .ZN(I38220) );
INV_X32 U_g29159 ( .A(I38220), .ZN(g29159) );
INV_X32 U_I38223 ( .A(g29106), .ZN(I38223) );
INV_X32 U_g29160 ( .A(I38223), .ZN(g29160) );
INV_X32 U_I38226 ( .A(g29108), .ZN(I38226) );
INV_X32 U_g29161 ( .A(I38226), .ZN(g29161) );
INV_X32 U_I38229 ( .A(g28950), .ZN(I38229) );
INV_X32 U_g29162 ( .A(I38229), .ZN(g29162) );
INV_X32 U_I38232 ( .A(g29117), .ZN(I38232) );
INV_X32 U_g29163 ( .A(I38232), .ZN(g29163) );
INV_X32 U_I38235 ( .A(g29118), .ZN(I38235) );
INV_X32 U_g29164 ( .A(I38235), .ZN(g29164) );
INV_X32 U_I38238 ( .A(g29119), .ZN(I38238) );
INV_X32 U_g29165 ( .A(I38238), .ZN(g29165) );
INV_X32 U_I38241 ( .A(g28832), .ZN(I38241) );
INV_X32 U_g29166 ( .A(I38241), .ZN(g29166) );
INV_X32 U_I38245 ( .A(g28920), .ZN(I38245) );
INV_X32 U_g29168 ( .A(I38245), .ZN(g29168) );
INV_X32 U_I38250 ( .A(g28941), .ZN(I38250) );
INV_X32 U_g29171 ( .A(I38250), .ZN(g29171) );
INV_X32 U_I38258 ( .A(g28963), .ZN(I38258) );
INV_X32 U_g29177 ( .A(I38258), .ZN(g29177) );
INV_X32 U_I38272 ( .A(g29013), .ZN(I38272) );
INV_X32 U_g29189 ( .A(I38272), .ZN(g29189) );
INV_X32 U_I38275 ( .A(g28987), .ZN(I38275) );
INV_X32 U_g29190 ( .A(I38275), .ZN(g29190) );
INV_X32 U_I38278 ( .A(g28963), .ZN(I38278) );
INV_X32 U_g29191 ( .A(I38278), .ZN(g29191) );
INV_X32 U_g29192 ( .A(g28954), .ZN(g29192) );
INV_X32 U_I38282 ( .A(g28941), .ZN(I38282) );
INV_X32 U_g29193 ( .A(I38282), .ZN(g29193) );
INV_X32 U_I38321 ( .A(g29113), .ZN(I38321) );
INV_X32 U_g29230 ( .A(I38321), .ZN(g29230) );
INV_X32 U_I38330 ( .A(g29120), .ZN(I38330) );
INV_X32 U_g29237 ( .A(I38330), .ZN(g29237) );
INV_X32 U_I38339 ( .A(g29120), .ZN(I38339) );
INV_X32 U_g29244 ( .A(I38339), .ZN(g29244) );
INV_X32 U_I38342 ( .A(g28886), .ZN(I38342) );
INV_X32 U_g29245 ( .A(I38342), .ZN(g29245) );
INV_X32 U_I38345 ( .A(g29109), .ZN(I38345) );
INV_X32 U_g29246 ( .A(I38345), .ZN(g29246) );
INV_X32 U_I38348 ( .A(g28874), .ZN(I38348) );
INV_X32 U_g29247 ( .A(I38348), .ZN(g29247) );
INV_X32 U_I38352 ( .A(g29110), .ZN(I38352) );
INV_X32 U_g29249 ( .A(I38352), .ZN(g29249) );
INV_X32 U_I38355 ( .A(g29039), .ZN(I38355) );
INV_X32 U_g29250 ( .A(I38355), .ZN(g29250) );
INV_X32 U_I38360 ( .A(g29111), .ZN(I38360) );
INV_X32 U_g29253 ( .A(I38360), .ZN(g29253) );
INV_X32 U_I38363 ( .A(g29016), .ZN(I38363) );
INV_X32 U_g29254 ( .A(I38363), .ZN(g29254) );
INV_X32 U_I38369 ( .A(g29112), .ZN(I38369) );
INV_X32 U_g29258 ( .A(I38369), .ZN(g29258) );
INV_X32 U_g29266 ( .A(g28741), .ZN(g29266) );
INV_X32 U_I38386 ( .A(g28734), .ZN(I38386) );
INV_X32 U_g29267 ( .A(I38386), .ZN(g29267) );
INV_X32 U_g29268 ( .A(g28751), .ZN(g29268) );
INV_X32 U_g29269 ( .A(g28755), .ZN(g29269) );
INV_X32 U_I38391 ( .A(g28730), .ZN(I38391) );
INV_X32 U_g29270 ( .A(I38391), .ZN(g29270) );
INV_X32 U_g29271 ( .A(g28764), .ZN(g29271) );
INV_X32 U_g29272 ( .A(g28768), .ZN(g29272) );
INV_X32 U_I38396 ( .A(g28727), .ZN(I38396) );
INV_X32 U_g29273 ( .A(I38396), .ZN(g29273) );
INV_X32 U_g29274 ( .A(g28775), .ZN(g29274) );
INV_X32 U_g29275 ( .A(g28779), .ZN(g29275) );
INV_X32 U_I38401 ( .A(g28725), .ZN(I38401) );
INV_X32 U_g29276 ( .A(I38401), .ZN(g29276) );
INV_X32 U_g29277 ( .A(g28785), .ZN(g29277) );
INV_X32 U_I38405 ( .A(g28723), .ZN(I38405) );
INV_X32 U_g29278 ( .A(I38405), .ZN(g29278) );
INV_X32 U_I38408 ( .A(g28721), .ZN(I38408) );
INV_X32 U_g29279 ( .A(I38408), .ZN(g29279) );
INV_X32 U_g29280 ( .A(g28791), .ZN(g29280) );
INV_X32 U_I38412 ( .A(g28720), .ZN(I38412) );
INV_X32 U_g29281 ( .A(I38412), .ZN(g29281) );
INV_X32 U_g29282 ( .A(g28796), .ZN(g29282) );
INV_X32 U_g29283 ( .A(g28799), .ZN(g29283) );
INV_X32 U_g29285 ( .A(g28804), .ZN(g29285) );
INV_X32 U_g29286 ( .A(g28807), .ZN(g29286) );
INV_X32 U_g29287 ( .A(g28810), .ZN(g29287) );
INV_X32 U_I38421 ( .A(g28740), .ZN(I38421) );
INV_X32 U_g29288 ( .A(I38421), .ZN(g29288) );
INV_X32 U_g29290 ( .A(g28814), .ZN(g29290) );
INV_X32 U_g29291 ( .A(g28817), .ZN(g29291) );
INV_X32 U_g29292 ( .A(g28820), .ZN(g29292) );
INV_X32 U_I38428 ( .A(g28732), .ZN(I38428) );
INV_X32 U_g29293 ( .A(I38428), .ZN(g29293) );
INV_X32 U_g29295 ( .A(g28823), .ZN(g29295) );
INV_X32 U_g29296 ( .A(g28826), .ZN(g29296) );
INV_X32 U_I38434 ( .A(g28735), .ZN(I38434) );
INV_X32 U_g29297 ( .A(I38434), .ZN(g29297) );
INV_X32 U_I38437 ( .A(g28736), .ZN(I38437) );
INV_X32 U_g29298 ( .A(I38437), .ZN(g29298) );
INV_X32 U_I38440 ( .A(g28738), .ZN(I38440) );
INV_X32 U_g29299 ( .A(I38440), .ZN(g29299) );
INV_X32 U_g29301 ( .A(g28829), .ZN(g29301) );
INV_X32 U_I38447 ( .A(g28744), .ZN(I38447) );
INV_X32 U_g29304 ( .A(I38447), .ZN(g29304) );
INV_X32 U_I38450 ( .A(g28745), .ZN(I38450) );
INV_X32 U_g29305 ( .A(I38450), .ZN(g29305) );
INV_X32 U_I38453 ( .A(g28746), .ZN(I38453) );
INV_X32 U_g29306 ( .A(I38453), .ZN(g29306) );
INV_X32 U_I38456 ( .A(g28747), .ZN(I38456) );
INV_X32 U_g29307 ( .A(I38456), .ZN(g29307) );
INV_X32 U_I38459 ( .A(g28749), .ZN(I38459) );
INV_X32 U_g29308 ( .A(I38459), .ZN(g29308) );
INV_X32 U_I38462 ( .A(g29120), .ZN(I38462) );
INV_X32 U_g29309 ( .A(I38462), .ZN(g29309) );
INV_X32 U_I38466 ( .A(g28754), .ZN(I38466) );
INV_X32 U_g29311 ( .A(I38466), .ZN(g29311) );
INV_X32 U_I38471 ( .A(g28758), .ZN(I38471) );
INV_X32 U_g29314 ( .A(I38471), .ZN(g29314) );
INV_X32 U_I38474 ( .A(g28759), .ZN(I38474) );
INV_X32 U_g29315 ( .A(I38474), .ZN(g29315) );
INV_X32 U_I38477 ( .A(g28760), .ZN(I38477) );
INV_X32 U_g29316 ( .A(I38477), .ZN(g29316) );
INV_X32 U_I38480 ( .A(g28761), .ZN(I38480) );
INV_X32 U_g29317 ( .A(I38480), .ZN(g29317) );
INV_X32 U_I38483 ( .A(g28990), .ZN(I38483) );
INV_X32 U_g29318 ( .A(I38483), .ZN(g29318) );
INV_X32 U_I38486 ( .A(g28763), .ZN(I38486) );
INV_X32 U_g29319 ( .A(I38486), .ZN(g29319) );
INV_X32 U_I38491 ( .A(g28767), .ZN(I38491) );
INV_X32 U_g29322 ( .A(I38491), .ZN(g29322) );
INV_X32 U_I38496 ( .A(g28771), .ZN(I38496) );
INV_X32 U_g29325 ( .A(I38496), .ZN(g29325) );
INV_X32 U_I38499 ( .A(g28772), .ZN(I38499) );
INV_X32 U_g29326 ( .A(I38499), .ZN(g29326) );
INV_X32 U_I38502 ( .A(g28773), .ZN(I38502) );
INV_X32 U_g29327 ( .A(I38502), .ZN(g29327) );
INV_X32 U_I38505 ( .A(g28774), .ZN(I38505) );
INV_X32 U_g29328 ( .A(I38505), .ZN(g29328) );
INV_X32 U_I38510 ( .A(g28778), .ZN(I38510) );
INV_X32 U_g29331 ( .A(I38510), .ZN(g29331) );
INV_X32 U_I38515 ( .A(g28782), .ZN(I38515) );
INV_X32 U_g29334 ( .A(I38515), .ZN(g29334) );
INV_X32 U_I38518 ( .A(g28783), .ZN(I38518) );
INV_X32 U_g29335 ( .A(I38518), .ZN(g29335) );
INV_X32 U_I38524 ( .A(g28788), .ZN(I38524) );
INV_X32 U_g29339 ( .A(I38524), .ZN(g29339) );
INV_X32 U_I38536 ( .A(g28920), .ZN(I38536) );
INV_X32 U_g29349 ( .A(I38536), .ZN(g29349) );
INV_X32 U_I38539 ( .A(g29113), .ZN(I38539) );
INV_X32 U_g29350 ( .A(I38539), .ZN(g29350) );
INV_X32 U_g29356 ( .A(g29120), .ZN(g29356) );
INV_X32 U_g29358 ( .A(g29120), .ZN(g29358) );
INV_X32 U_I38548 ( .A(g28903), .ZN(I38548) );
INV_X32 U_g29359 ( .A(I38548), .ZN(g29359) );
INV_X32 U_g29360 ( .A(g28871), .ZN(g29360) );
INV_X32 U_g29361 ( .A(g28877), .ZN(g29361) );
INV_X32 U_g29362 ( .A(g28883), .ZN(g29362) );
INV_X32 U_g29363 ( .A(g28889), .ZN(g29363) );
INV_X32 U_g29364 ( .A(g28894), .ZN(g29364) );
INV_X32 U_g29365 ( .A(g28900), .ZN(g29365) );
INV_X32 U_g29366 ( .A(g28906), .ZN(g29366) );
INV_X32 U_g29367 ( .A(g28911), .ZN(g29367) );
INV_X32 U_g29368 ( .A(g28916), .ZN(g29368) );
INV_X32 U_g29369 ( .A(g28925), .ZN(g29369) );
INV_X32 U_g29370 ( .A(g28928), .ZN(g29370) );
INV_X32 U_g29371 ( .A(g28932), .ZN(g29371) );
INV_X32 U_g29372 ( .A(g28937), .ZN(g29372) );
INV_X32 U_g29373 ( .A(g28945), .ZN(g29373) );
INV_X32 U_g29374 ( .A(g28951), .ZN(g29374) );
INV_X32 U_g29375 ( .A(g28955), .ZN(g29375) );
INV_X32 U_g29376 ( .A(g28959), .ZN(g29376) );
INV_X32 U_g29377 ( .A(g28967), .ZN(g29377) );
INV_X32 U_g29378 ( .A(g28972), .ZN(g29378) );
INV_X32 U_g29379 ( .A(g28975), .ZN(g29379) );
INV_X32 U_g29380 ( .A(g28979), .ZN(g29380) );
INV_X32 U_g29381 ( .A(g28983), .ZN(g29381) );
INV_X32 U_g29382 ( .A(g28993), .ZN(g29382) );
INV_X32 U_g29383 ( .A(g28998), .ZN(g29383) );
INV_X32 U_g29384 ( .A(g29002), .ZN(g29384) );
INV_X32 U_g29385 ( .A(g29005), .ZN(g29385) );
INV_X32 U_g29386 ( .A(g29010), .ZN(g29386) );
INV_X32 U_g29387 ( .A(g29019), .ZN(g29387) );
INV_X32 U_g29388 ( .A(g29023), .ZN(g29388) );
INV_X32 U_g29389 ( .A(g29027), .ZN(g29389) );
INV_X32 U_g29390 ( .A(g29032), .ZN(g29390) );
INV_X32 U_g29391 ( .A(g29035), .ZN(g29391) );
INV_X32 U_g29392 ( .A(g29042), .ZN(g29392) );
INV_X32 U_g29393 ( .A(g29046), .ZN(g29393) );
INV_X32 U_g29394 ( .A(g29050), .ZN(g29394) );
INV_X32 U_g29395 ( .A(g29054), .ZN(g29395) );
INV_X32 U_g29396 ( .A(g29057), .ZN(g29396) );
INV_X32 U_g29397 ( .A(g29065), .ZN(g29397) );
INV_X32 U_g29398 ( .A(g29069), .ZN(g29398) );
INV_X32 U_I38591 ( .A(g28987), .ZN(I38591) );
INV_X32 U_g29400 ( .A(I38591), .ZN(g29400) );
INV_X32 U_I38594 ( .A(g28990), .ZN(I38594) );
INV_X32 U_g29401 ( .A(I38594), .ZN(g29401) );
INV_X32 U_g29402 ( .A(g29077), .ZN(g29402) );
INV_X32 U_I38599 ( .A(g29013), .ZN(I38599) );
INV_X32 U_g29404 ( .A(I38599), .ZN(g29404) );
INV_X32 U_I38602 ( .A(g29016), .ZN(I38602) );
INV_X32 U_g29405 ( .A(I38602), .ZN(g29405) );
INV_X32 U_I38606 ( .A(g29039), .ZN(I38606) );
INV_X32 U_g29407 ( .A(I38606), .ZN(g29407) );
INV_X32 U_I38609 ( .A(g28874), .ZN(I38609) );
INV_X32 U_g29408 ( .A(I38609), .ZN(g29408) );
INV_X32 U_I38613 ( .A(g28886), .ZN(I38613) );
INV_X32 U_g29410 ( .A(I38613), .ZN(g29410) );
INV_X32 U_I38617 ( .A(g28903), .ZN(I38617) );
INV_X32 U_g29412 ( .A(I38617), .ZN(g29412) );
INV_X32 U_I38620 ( .A(g29246), .ZN(I38620) );
INV_X32 U_g29413 ( .A(I38620), .ZN(g29413) );
INV_X32 U_I38623 ( .A(g29293), .ZN(I38623) );
INV_X32 U_g29414 ( .A(I38623), .ZN(g29414) );
INV_X32 U_I38626 ( .A(g29297), .ZN(I38626) );
INV_X32 U_g29415 ( .A(I38626), .ZN(g29415) );
INV_X32 U_I38629 ( .A(g29304), .ZN(I38629) );
INV_X32 U_g29416 ( .A(I38629), .ZN(g29416) );
INV_X32 U_I38632 ( .A(g29298), .ZN(I38632) );
INV_X32 U_g29417 ( .A(I38632), .ZN(g29417) );
INV_X32 U_I38635 ( .A(g29305), .ZN(I38635) );
INV_X32 U_g29418 ( .A(I38635), .ZN(g29418) );
INV_X32 U_I38638 ( .A(g29311), .ZN(I38638) );
INV_X32 U_g29419 ( .A(I38638), .ZN(g29419) );
INV_X32 U_I38641 ( .A(g29249), .ZN(I38641) );
INV_X32 U_g29420 ( .A(I38641), .ZN(g29420) );
INV_X32 U_I38644 ( .A(g29299), .ZN(I38644) );
INV_X32 U_g29421 ( .A(I38644), .ZN(g29421) );
INV_X32 U_I38647 ( .A(g29306), .ZN(I38647) );
INV_X32 U_g29422 ( .A(I38647), .ZN(g29422) );
INV_X32 U_I38650 ( .A(g29314), .ZN(I38650) );
INV_X32 U_g29423 ( .A(I38650), .ZN(g29423) );
INV_X32 U_I38653 ( .A(g29307), .ZN(I38653) );
INV_X32 U_g29424 ( .A(I38653), .ZN(g29424) );
INV_X32 U_I38656 ( .A(g29315), .ZN(I38656) );
INV_X32 U_g29425 ( .A(I38656), .ZN(g29425) );
INV_X32 U_I38659 ( .A(g29322), .ZN(I38659) );
INV_X32 U_g29426 ( .A(I38659), .ZN(g29426) );
INV_X32 U_I38662 ( .A(g29253), .ZN(I38662) );
INV_X32 U_g29427 ( .A(I38662), .ZN(g29427) );
INV_X32 U_I38665 ( .A(g29412), .ZN(I38665) );
INV_X32 U_g29428 ( .A(I38665), .ZN(g29428) );
INV_X32 U_I38668 ( .A(g29168), .ZN(I38668) );
INV_X32 U_g29429 ( .A(I38668), .ZN(g29429) );
INV_X32 U_I38671 ( .A(g29171), .ZN(I38671) );
INV_X32 U_g29430 ( .A(I38671), .ZN(g29430) );
INV_X32 U_I38674 ( .A(g29177), .ZN(I38674) );
INV_X32 U_g29431 ( .A(I38674), .ZN(g29431) );
INV_X32 U_I38677 ( .A(g29400), .ZN(I38677) );
INV_X32 U_g29432 ( .A(I38677), .ZN(g29432) );
INV_X32 U_I38680 ( .A(g29404), .ZN(I38680) );
INV_X32 U_g29433 ( .A(I38680), .ZN(g29433) );
INV_X32 U_I38683 ( .A(g29308), .ZN(I38683) );
INV_X32 U_g29434 ( .A(I38683), .ZN(g29434) );
INV_X32 U_I38686 ( .A(g29316), .ZN(I38686) );
INV_X32 U_g29435 ( .A(I38686), .ZN(g29435) );
INV_X32 U_I38689 ( .A(g29325), .ZN(I38689) );
INV_X32 U_g29436 ( .A(I38689), .ZN(g29436) );
INV_X32 U_I38692 ( .A(g29317), .ZN(I38692) );
INV_X32 U_g29437 ( .A(I38692), .ZN(g29437) );
INV_X32 U_I38695 ( .A(g29326), .ZN(I38695) );
INV_X32 U_g29438 ( .A(I38695), .ZN(g29438) );
INV_X32 U_I38698 ( .A(g29331), .ZN(I38698) );
INV_X32 U_g29439 ( .A(I38698), .ZN(g29439) );
INV_X32 U_I38701 ( .A(g29401), .ZN(I38701) );
INV_X32 U_g29440 ( .A(I38701), .ZN(g29440) );
INV_X32 U_I38704 ( .A(g29405), .ZN(I38704) );
INV_X32 U_g29441 ( .A(I38704), .ZN(g29441) );
INV_X32 U_I38707 ( .A(g29407), .ZN(I38707) );
INV_X32 U_g29442 ( .A(I38707), .ZN(g29442) );
INV_X32 U_I38710 ( .A(g29408), .ZN(I38710) );
INV_X32 U_g29443 ( .A(I38710), .ZN(g29443) );
INV_X32 U_I38713 ( .A(g29410), .ZN(I38713) );
INV_X32 U_g29444 ( .A(I38713), .ZN(g29444) );
INV_X32 U_I38716 ( .A(g29230), .ZN(I38716) );
INV_X32 U_g29445 ( .A(I38716), .ZN(g29445) );
INV_X32 U_I38719 ( .A(g29258), .ZN(I38719) );
INV_X32 U_g29446 ( .A(I38719), .ZN(g29446) );
INV_X32 U_I38722 ( .A(g29319), .ZN(I38722) );
INV_X32 U_g29447 ( .A(I38722), .ZN(g29447) );
INV_X32 U_I38725 ( .A(g29327), .ZN(I38725) );
INV_X32 U_g29448 ( .A(I38725), .ZN(g29448) );
INV_X32 U_I38728 ( .A(g29334), .ZN(I38728) );
INV_X32 U_g29449 ( .A(I38728), .ZN(g29449) );
INV_X32 U_I38731 ( .A(g29328), .ZN(I38731) );
INV_X32 U_g29450 ( .A(I38731), .ZN(g29450) );
INV_X32 U_I38734 ( .A(g29335), .ZN(I38734) );
INV_X32 U_g29451 ( .A(I38734), .ZN(g29451) );
INV_X32 U_I38737 ( .A(g29339), .ZN(I38737) );
INV_X32 U_g29452 ( .A(I38737), .ZN(g29452) );
INV_X32 U_I38740 ( .A(g29288), .ZN(I38740) );
INV_X32 U_g29453 ( .A(I38740), .ZN(g29453) );
INV_X32 U_I38743 ( .A(g29267), .ZN(I38743) );
INV_X32 U_g29454 ( .A(I38743), .ZN(g29454) );
INV_X32 U_I38746 ( .A(g29270), .ZN(I38746) );
INV_X32 U_g29455 ( .A(I38746), .ZN(g29455) );
INV_X32 U_I38749 ( .A(g29273), .ZN(I38749) );
INV_X32 U_g29456 ( .A(I38749), .ZN(g29456) );
INV_X32 U_I38752 ( .A(g29276), .ZN(I38752) );
INV_X32 U_g29457 ( .A(I38752), .ZN(g29457) );
INV_X32 U_I38755 ( .A(g29278), .ZN(I38755) );
INV_X32 U_g29458 ( .A(I38755), .ZN(g29458) );
INV_X32 U_I38758 ( .A(g29279), .ZN(I38758) );
INV_X32 U_g29459 ( .A(I38758), .ZN(g29459) );
INV_X32 U_I38761 ( .A(g29281), .ZN(I38761) );
INV_X32 U_g29460 ( .A(I38761), .ZN(g29460) );
INV_X32 U_I38764 ( .A(g29237), .ZN(I38764) );
INV_X32 U_g29461 ( .A(I38764), .ZN(g29461) );
INV_X32 U_I38767 ( .A(g29244), .ZN(I38767) );
INV_X32 U_g29462 ( .A(I38767), .ZN(g29462) );
INV_X32 U_I38770 ( .A(g29309), .ZN(I38770) );
INV_X32 U_g29463 ( .A(I38770), .ZN(g29463) );
INV_X32 U_g29491 ( .A(g29350), .ZN(g29491) );
INV_X32 U_I38801 ( .A(g29358), .ZN(I38801) );
INV_X32 U_g29495 ( .A(I38801), .ZN(g29495) );
INV_X32 U_I38804 ( .A(g29353), .ZN(I38804) );
INV_X32 U_g29496 ( .A(I38804), .ZN(g29496) );
INV_X32 U_I38807 ( .A(g29356), .ZN(I38807) );
INV_X32 U_g29497 ( .A(I38807), .ZN(g29497) );
INV_X32 U_I38817 ( .A(g29354), .ZN(I38817) );
INV_X32 U_g29499 ( .A(I38817), .ZN(g29499) );
INV_X32 U_I38827 ( .A(g29355), .ZN(I38827) );
INV_X32 U_g29501 ( .A(I38827), .ZN(g29501) );
INV_X32 U_I38838 ( .A(g29357), .ZN(I38838) );
INV_X32 U_g29504 ( .A(I38838), .ZN(g29504) );
INV_X32 U_I38848 ( .A(g29167), .ZN(I38848) );
INV_X32 U_g29506 ( .A(I38848), .ZN(g29506) );
INV_X32 U_I38851 ( .A(g29169), .ZN(I38851) );
INV_X32 U_g29507 ( .A(I38851), .ZN(g29507) );
INV_X32 U_I38854 ( .A(g29170), .ZN(I38854) );
INV_X32 U_g29508 ( .A(I38854), .ZN(g29508) );
INV_X32 U_I38857 ( .A(g29172), .ZN(I38857) );
INV_X32 U_g29509 ( .A(I38857), .ZN(g29509) );
INV_X32 U_I38860 ( .A(g29173), .ZN(I38860) );
INV_X32 U_g29510 ( .A(I38860), .ZN(g29510) );
INV_X32 U_I38863 ( .A(g29178), .ZN(I38863) );
INV_X32 U_g29511 ( .A(I38863), .ZN(g29511) );
INV_X32 U_I38866 ( .A(g29179), .ZN(I38866) );
INV_X32 U_g29512 ( .A(I38866), .ZN(g29512) );
INV_X32 U_I38869 ( .A(g29181), .ZN(I38869) );
INV_X32 U_g29513 ( .A(I38869), .ZN(g29513) );
INV_X32 U_I38872 ( .A(g29182), .ZN(I38872) );
INV_X32 U_g29514 ( .A(I38872), .ZN(g29514) );
INV_X32 U_I38875 ( .A(g29184), .ZN(I38875) );
INV_X32 U_g29515 ( .A(I38875), .ZN(g29515) );
INV_X32 U_I38878 ( .A(g29185), .ZN(I38878) );
INV_X32 U_g29516 ( .A(I38878), .ZN(g29516) );
INV_X32 U_I38881 ( .A(g29187), .ZN(I38881) );
INV_X32 U_g29517 ( .A(I38881), .ZN(g29517) );
INV_X32 U_I38885 ( .A(g29192), .ZN(I38885) );
INV_X32 U_g29519 ( .A(I38885), .ZN(g29519) );
INV_X32 U_I38898 ( .A(g29194), .ZN(I38898) );
INV_X32 U_g29530 ( .A(I38898), .ZN(g29530) );
INV_X32 U_I38905 ( .A(g29197), .ZN(I38905) );
INV_X32 U_g29535 ( .A(I38905), .ZN(g29535) );
INV_X32 U_I38909 ( .A(g29198), .ZN(I38909) );
INV_X32 U_g29537 ( .A(I38909), .ZN(g29537) );
INV_X32 U_I38916 ( .A(g29201), .ZN(I38916) );
INV_X32 U_g29542 ( .A(I38916), .ZN(g29542) );
INV_X32 U_I38920 ( .A(g29204), .ZN(I38920) );
INV_X32 U_g29544 ( .A(I38920), .ZN(g29544) );
INV_X32 U_I38924 ( .A(g29205), .ZN(I38924) );
INV_X32 U_g29546 ( .A(I38924), .ZN(g29546) );
INV_X32 U_I38931 ( .A(g29209), .ZN(I38931) );
INV_X32 U_g29551 ( .A(I38931), .ZN(g29551) );
INV_X32 U_I38936 ( .A(g29212), .ZN(I38936) );
INV_X32 U_g29554 ( .A(I38936), .ZN(g29554) );
INV_X32 U_I38940 ( .A(g29213), .ZN(I38940) );
INV_X32 U_g29556 ( .A(I38940), .ZN(g29556) );
INV_X32 U_I38947 ( .A(g29218), .ZN(I38947) );
INV_X32 U_g29561 ( .A(I38947), .ZN(g29561) );
INV_X32 U_I38951 ( .A(g29221), .ZN(I38951) );
INV_X32 U_g29563 ( .A(I38951), .ZN(g29563) );
INV_X32 U_I38958 ( .A(g29226), .ZN(I38958) );
INV_X32 U_g29568 ( .A(I38958), .ZN(g29568) );
INV_X32 U_I38975 ( .A(g29348), .ZN(I38975) );
INV_X32 U_g29583 ( .A(I38975), .ZN(g29583) );
INV_X32 U_I38999 ( .A(g29496), .ZN(I38999) );
INV_X32 U_g29627 ( .A(I38999), .ZN(g29627) );
INV_X32 U_I39002 ( .A(g29506), .ZN(I39002) );
INV_X32 U_g29628 ( .A(I39002), .ZN(g29628) );
INV_X32 U_I39005 ( .A(g29507), .ZN(I39005) );
INV_X32 U_g29629 ( .A(I39005), .ZN(g29629) );
INV_X32 U_I39008 ( .A(g29509), .ZN(I39008) );
INV_X32 U_g29630 ( .A(I39008), .ZN(g29630) );
INV_X32 U_I39011 ( .A(g29530), .ZN(I39011) );
INV_X32 U_g29631 ( .A(I39011), .ZN(g29631) );
INV_X32 U_I39014 ( .A(g29535), .ZN(I39014) );
INV_X32 U_g29632 ( .A(I39014), .ZN(g29632) );
INV_X32 U_I39017 ( .A(g29542), .ZN(I39017) );
INV_X32 U_g29633 ( .A(I39017), .ZN(g29633) );
INV_X32 U_I39020 ( .A(g29499), .ZN(I39020) );
INV_X32 U_g29634 ( .A(I39020), .ZN(g29634) );
INV_X32 U_I39023 ( .A(g29508), .ZN(I39023) );
INV_X32 U_g29635 ( .A(I39023), .ZN(g29635) );
INV_X32 U_I39026 ( .A(g29510), .ZN(I39026) );
INV_X32 U_g29636 ( .A(I39026), .ZN(g29636) );
INV_X32 U_I39029 ( .A(g29512), .ZN(I39029) );
INV_X32 U_g29637 ( .A(I39029), .ZN(g29637) );
INV_X32 U_I39032 ( .A(g29537), .ZN(I39032) );
INV_X32 U_g29638 ( .A(I39032), .ZN(g29638) );
INV_X32 U_I39035 ( .A(g29544), .ZN(I39035) );
INV_X32 U_g29639 ( .A(I39035), .ZN(g29639) );
INV_X32 U_I39038 ( .A(g29551), .ZN(I39038) );
INV_X32 U_g29640 ( .A(I39038), .ZN(g29640) );
INV_X32 U_I39041 ( .A(g29501), .ZN(I39041) );
INV_X32 U_g29641 ( .A(I39041), .ZN(g29641) );
INV_X32 U_I39044 ( .A(g29511), .ZN(I39044) );
INV_X32 U_g29642 ( .A(I39044), .ZN(g29642) );
INV_X32 U_I39047 ( .A(g29513), .ZN(I39047) );
INV_X32 U_g29643 ( .A(I39047), .ZN(g29643) );
INV_X32 U_I39050 ( .A(g29515), .ZN(I39050) );
INV_X32 U_g29644 ( .A(I39050), .ZN(g29644) );
INV_X32 U_I39053 ( .A(g29546), .ZN(I39053) );
INV_X32 U_g29645 ( .A(I39053), .ZN(g29645) );
INV_X32 U_I39056 ( .A(g29554), .ZN(I39056) );
INV_X32 U_g29646 ( .A(I39056), .ZN(g29646) );
INV_X32 U_I39059 ( .A(g29561), .ZN(I39059) );
INV_X32 U_g29647 ( .A(I39059), .ZN(g29647) );
INV_X32 U_I39062 ( .A(g29504), .ZN(I39062) );
INV_X32 U_g29648 ( .A(I39062), .ZN(g29648) );
INV_X32 U_I39065 ( .A(g29514), .ZN(I39065) );
INV_X32 U_g29649 ( .A(I39065), .ZN(g29649) );
INV_X32 U_I39068 ( .A(g29516), .ZN(I39068) );
INV_X32 U_g29650 ( .A(I39068), .ZN(g29650) );
INV_X32 U_I39071 ( .A(g29517), .ZN(I39071) );
INV_X32 U_g29651 ( .A(I39071), .ZN(g29651) );
INV_X32 U_I39074 ( .A(g29556), .ZN(I39074) );
INV_X32 U_g29652 ( .A(I39074), .ZN(g29652) );
INV_X32 U_I39077 ( .A(g29563), .ZN(I39077) );
INV_X32 U_g29653 ( .A(I39077), .ZN(g29653) );
INV_X32 U_I39080 ( .A(g29568), .ZN(I39080) );
INV_X32 U_g29654 ( .A(I39080), .ZN(g29654) );
INV_X32 U_I39083 ( .A(g29519), .ZN(I39083) );
INV_X32 U_g29655 ( .A(I39083), .ZN(g29655) );
INV_X32 U_I39086 ( .A(g29497), .ZN(I39086) );
INV_X32 U_g29656 ( .A(I39086), .ZN(g29656) );
INV_X32 U_I39089 ( .A(g29495), .ZN(I39089) );
INV_X32 U_g29657 ( .A(I39089), .ZN(g29657) );
INV_X32 U_g29658 ( .A(g29574), .ZN(g29658) );
INV_X32 U_g29659 ( .A(g29571), .ZN(g29659) );
INV_X32 U_g29660 ( .A(g29578), .ZN(g29660) );
INV_X32 U_g29661 ( .A(g29576), .ZN(g29661) );
INV_X32 U_g29662 ( .A(g29570), .ZN(g29662) );
INV_X32 U_g29664 ( .A(g29552), .ZN(g29664) );
INV_X32 U_g29666 ( .A(g29577), .ZN(g29666) );
INV_X32 U_g29668 ( .A(g29569), .ZN(g29668) );
INV_X32 U_g29673 ( .A(g29583), .ZN(g29673) );
INV_X32 U_I39121 ( .A(g29579), .ZN(I39121) );
INV_X32 U_g29689 ( .A(I39121), .ZN(g29689) );
INV_X32 U_I39124 ( .A(g29606), .ZN(I39124) );
INV_X32 U_g29690 ( .A(I39124), .ZN(g29690) );
INV_X32 U_I39127 ( .A(g29608), .ZN(I39127) );
INV_X32 U_g29691 ( .A(I39127), .ZN(g29691) );
INV_X32 U_I39130 ( .A(g29580), .ZN(I39130) );
INV_X32 U_g29692 ( .A(I39130), .ZN(g29692) );
INV_X32 U_I39133 ( .A(g29609), .ZN(I39133) );
INV_X32 U_g29693 ( .A(I39133), .ZN(g29693) );
INV_X32 U_I39136 ( .A(g29611), .ZN(I39136) );
INV_X32 U_g29694 ( .A(I39136), .ZN(g29694) );
INV_X32 U_I39139 ( .A(g29612), .ZN(I39139) );
INV_X32 U_g29695 ( .A(I39139), .ZN(g29695) );
INV_X32 U_I39142 ( .A(g29581), .ZN(I39142) );
INV_X32 U_g29696 ( .A(I39142), .ZN(g29696) );
INV_X32 U_I39145 ( .A(g29613), .ZN(I39145) );
INV_X32 U_g29697 ( .A(I39145), .ZN(g29697) );
INV_X32 U_I39148 ( .A(g29616), .ZN(I39148) );
INV_X32 U_g29698 ( .A(I39148), .ZN(g29698) );
INV_X32 U_I39151 ( .A(g29617), .ZN(I39151) );
INV_X32 U_g29699 ( .A(I39151), .ZN(g29699) );
INV_X32 U_I39154 ( .A(g29582), .ZN(I39154) );
INV_X32 U_g29700 ( .A(I39154), .ZN(g29700) );
INV_X32 U_I39157 ( .A(g29618), .ZN(I39157) );
INV_X32 U_g29701 ( .A(I39157), .ZN(g29701) );
INV_X32 U_I39160 ( .A(g29620), .ZN(I39160) );
INV_X32 U_g29702 ( .A(I39160), .ZN(g29702) );
INV_X32 U_I39164 ( .A(g29621), .ZN(I39164) );
INV_X32 U_g29704 ( .A(I39164), .ZN(g29704) );
INV_X32 U_I39168 ( .A(g29623), .ZN(I39168) );
INV_X32 U_g29708 ( .A(I39168), .ZN(g29708) );
INV_X32 U_g29716 ( .A(g29498), .ZN(g29716) );
INV_X32 U_g29724 ( .A(g29500), .ZN(g29724) );
INV_X32 U_g29726 ( .A(g29503), .ZN(g29726) );
INV_X32 U_g29739 ( .A(g29505), .ZN(g29739) );
INV_X32 U_I39234 ( .A(g29689), .ZN(I39234) );
INV_X32 U_g29794 ( .A(I39234), .ZN(g29794) );
INV_X32 U_I39237 ( .A(g29690), .ZN(I39237) );
INV_X32 U_g29795 ( .A(I39237), .ZN(g29795) );
INV_X32 U_I39240 ( .A(g29691), .ZN(I39240) );
INV_X32 U_g29796 ( .A(I39240), .ZN(g29796) );
INV_X32 U_I39243 ( .A(g29694), .ZN(I39243) );
INV_X32 U_g29797 ( .A(I39243), .ZN(g29797) );
INV_X32 U_I39246 ( .A(g29692), .ZN(I39246) );
INV_X32 U_g29798 ( .A(I39246), .ZN(g29798) );
INV_X32 U_I39249 ( .A(g29693), .ZN(I39249) );
INV_X32 U_g29799 ( .A(I39249), .ZN(g29799) );
INV_X32 U_I39252 ( .A(g29695), .ZN(I39252) );
INV_X32 U_g29800 ( .A(I39252), .ZN(g29800) );
INV_X32 U_I39255 ( .A(g29698), .ZN(I39255) );
INV_X32 U_g29801 ( .A(I39255), .ZN(g29801) );
INV_X32 U_I39258 ( .A(g29696), .ZN(I39258) );
INV_X32 U_g29802 ( .A(I39258), .ZN(g29802) );
INV_X32 U_I39261 ( .A(g29697), .ZN(I39261) );
INV_X32 U_g29803 ( .A(I39261), .ZN(g29803) );
INV_X32 U_I39264 ( .A(g29699), .ZN(I39264) );
INV_X32 U_g29804 ( .A(I39264), .ZN(g29804) );
INV_X32 U_I39267 ( .A(g29702), .ZN(I39267) );
INV_X32 U_g29805 ( .A(I39267), .ZN(g29805) );
INV_X32 U_I39270 ( .A(g29700), .ZN(I39270) );
INV_X32 U_g29806 ( .A(I39270), .ZN(g29806) );
INV_X32 U_I39273 ( .A(g29701), .ZN(I39273) );
INV_X32 U_g29807 ( .A(I39273), .ZN(g29807) );
INV_X32 U_I39276 ( .A(g29704), .ZN(I39276) );
INV_X32 U_g29808 ( .A(I39276), .ZN(g29808) );
INV_X32 U_I39279 ( .A(g29708), .ZN(I39279) );
INV_X32 U_g29809 ( .A(I39279), .ZN(g29809) );
INV_X32 U_g29823 ( .A(g29663), .ZN(g29823) );
INV_X32 U_g29829 ( .A(g29665), .ZN(g29829) );
INV_X32 U_g29835 ( .A(g29667), .ZN(g29835) );
INV_X32 U_g29840 ( .A(g29669), .ZN(g29840) );
INV_X32 U_g29844 ( .A(g29670), .ZN(g29844) );
INV_X32 U_g29848 ( .A(g29761), .ZN(g29848) );
INV_X32 U_g29849 ( .A(g29671), .ZN(g29849) );
INV_X32 U_g29853 ( .A(g29672), .ZN(g29853) );
INV_X32 U_g29857 ( .A(g29676), .ZN(g29857) );
INV_X32 U_g29861 ( .A(g29677), .ZN(g29861) );
INV_X32 U_g29865 ( .A(g29678), .ZN(g29865) );
INV_X32 U_g29869 ( .A(g29679), .ZN(g29869) );
INV_X32 U_g29873 ( .A(g29680), .ZN(g29873) );
INV_X32 U_g29877 ( .A(g29681), .ZN(g29877) );
INV_X32 U_g29881 ( .A(g29682), .ZN(g29881) );
INV_X32 U_g29885 ( .A(g29683), .ZN(g29885) );
INV_X32 U_g29889 ( .A(g29684), .ZN(g29889) );
INV_X32 U_g29893 ( .A(g29685), .ZN(g29893) );
INV_X32 U_g29897 ( .A(g29686), .ZN(g29897) );
INV_X32 U_g29901 ( .A(g29687), .ZN(g29901) );
INV_X32 U_g29905 ( .A(g29688), .ZN(g29905) );
INV_X32 U_I39398 ( .A(g29664), .ZN(I39398) );
INV_X32 U_g29932 ( .A(I39398), .ZN(g29932) );
INV_X32 U_I39401 ( .A(g29662), .ZN(I39401) );
INV_X32 U_g29933 ( .A(I39401), .ZN(g29933) );
INV_X32 U_I39404 ( .A(g29661), .ZN(I39404) );
INV_X32 U_g29934 ( .A(I39404), .ZN(g29934) );
INV_X32 U_I39407 ( .A(g29660), .ZN(I39407) );
INV_X32 U_g29935 ( .A(I39407), .ZN(g29935) );
INV_X32 U_I39411 ( .A(g29659), .ZN(I39411) );
INV_X32 U_g29937 ( .A(I39411), .ZN(g29937) );
INV_X32 U_I39414 ( .A(g29658), .ZN(I39414) );
INV_X32 U_g29938 ( .A(I39414), .ZN(g29938) );
INV_X32 U_I39418 ( .A(g29668), .ZN(I39418) );
INV_X32 U_g29940 ( .A(I39418), .ZN(g29940) );
INV_X32 U_I39423 ( .A(g29666), .ZN(I39423) );
INV_X32 U_g29943 ( .A(I39423), .ZN(g29943) );
INV_X32 U_I39454 ( .A(g29940), .ZN(I39454) );
INV_X32 U_g29972 ( .A(I39454), .ZN(g29972) );
INV_X32 U_I39457 ( .A(g29943), .ZN(I39457) );
INV_X32 U_g29973 ( .A(I39457), .ZN(g29973) );
INV_X32 U_I39460 ( .A(g29932), .ZN(I39460) );
INV_X32 U_g29974 ( .A(I39460), .ZN(g29974) );
INV_X32 U_I39463 ( .A(g29933), .ZN(I39463) );
INV_X32 U_g29975 ( .A(I39463), .ZN(g29975) );
INV_X32 U_I39466 ( .A(g29934), .ZN(I39466) );
INV_X32 U_g29976 ( .A(I39466), .ZN(g29976) );
INV_X32 U_I39469 ( .A(g29935), .ZN(I39469) );
INV_X32 U_g29977 ( .A(I39469), .ZN(g29977) );
INV_X32 U_I39472 ( .A(g29937), .ZN(I39472) );
INV_X32 U_g29978 ( .A(I39472), .ZN(g29978) );
INV_X32 U_I39475 ( .A(g29938), .ZN(I39475) );
INV_X32 U_g29979 ( .A(I39475), .ZN(g29979) );
INV_X32 U_g30036 ( .A(g29912), .ZN(g30036) );
INV_X32 U_g30040 ( .A(g29914), .ZN(g30040) );
INV_X32 U_g30044 ( .A(g29916), .ZN(g30044) );
INV_X32 U_g30048 ( .A(g29920), .ZN(g30048) );
INV_X32 U_I39550 ( .A(g29848), .ZN(I39550) );
INV_X32 U_g30052 ( .A(I39550), .ZN(g30052) );
INV_X32 U_I39573 ( .A(g29936), .ZN(I39573) );
INV_X32 U_g30076 ( .A(I39573), .ZN(g30076) );
INV_X32 U_I39577 ( .A(g29939), .ZN(I39577) );
INV_X32 U_g30078 ( .A(I39577), .ZN(g30078) );
INV_X32 U_I39585 ( .A(g29941), .ZN(I39585) );
INV_X32 U_g30084 ( .A(I39585), .ZN(g30084) );
INV_X32 U_I39622 ( .A(g30052), .ZN(I39622) );
INV_X32 U_g30119 ( .A(I39622), .ZN(g30119) );
INV_X32 U_I39625 ( .A(g30076), .ZN(I39625) );
INV_X32 U_g30120 ( .A(I39625), .ZN(g30120) );
INV_X32 U_I39628 ( .A(g30078), .ZN(I39628) );
INV_X32 U_g30121 ( .A(I39628), .ZN(g30121) );
INV_X32 U_I39631 ( .A(g30084), .ZN(I39631) );
INV_X32 U_g30122 ( .A(I39631), .ZN(g30122) );
INV_X32 U_I39635 ( .A(g30055), .ZN(I39635) );
INV_X32 U_g30124 ( .A(I39635), .ZN(g30124) );
INV_X32 U_I39638 ( .A(g30056), .ZN(I39638) );
INV_X32 U_g30125 ( .A(I39638), .ZN(g30125) );
INV_X32 U_I39641 ( .A(g30057), .ZN(I39641) );
INV_X32 U_g30126 ( .A(I39641), .ZN(g30126) );
INV_X32 U_I39647 ( .A(g30058), .ZN(I39647) );
INV_X32 U_g30130 ( .A(I39647), .ZN(g30130) );
INV_X32 U_g30134 ( .A(g30010), .ZN(g30134) );
INV_X32 U_g30139 ( .A(g30011), .ZN(g30139) );
INV_X32 U_g30143 ( .A(g30012), .ZN(g30143) );
INV_X32 U_g30147 ( .A(g30013), .ZN(g30147) );
INV_X32 U_g30151 ( .A(g30014), .ZN(g30151) );
INV_X32 U_g30155 ( .A(g30015), .ZN(g30155) );
INV_X32 U_g30159 ( .A(g30016), .ZN(g30159) );
INV_X32 U_g30163 ( .A(g30017), .ZN(g30163) );
INV_X32 U_g30167 ( .A(g30018), .ZN(g30167) );
INV_X32 U_g30171 ( .A(g30019), .ZN(g30171) );
INV_X32 U_g30175 ( .A(g30020), .ZN(g30175) );
INV_X32 U_g30179 ( .A(g30021), .ZN(g30179) );
INV_X32 U_g30183 ( .A(g30022), .ZN(g30183) );
INV_X32 U_g30187 ( .A(g30023), .ZN(g30187) );
INV_X32 U_g30191 ( .A(g30024), .ZN(g30191) );
INV_X32 U_g30195 ( .A(g30025), .ZN(g30195) );
INV_X32 U_g30199 ( .A(g30026), .ZN(g30199) );
INV_X32 U_g30203 ( .A(g30027), .ZN(g30203) );
INV_X32 U_g30207 ( .A(g30028), .ZN(g30207) );
INV_X32 U_g30211 ( .A(g30029), .ZN(g30211) );
INV_X32 U_I39674 ( .A(g30072), .ZN(I39674) );
INV_X32 U_g30215 ( .A(I39674), .ZN(g30215) );
INV_X32 U_g30229 ( .A(g30030), .ZN(g30229) );
INV_X32 U_g30233 ( .A(g30031), .ZN(g30233) );
INV_X32 U_g30237 ( .A(g30032), .ZN(g30237) );
INV_X32 U_g30241 ( .A(g30033), .ZN(g30241) );
INV_X32 U_I39761 ( .A(g30072), .ZN(I39761) );
INV_X32 U_g30306 ( .A(I39761), .ZN(g30306) );
INV_X32 U_I39764 ( .A(g30060), .ZN(I39764) );
INV_X32 U_g30307 ( .A(I39764), .ZN(g30307) );
INV_X32 U_I39767 ( .A(g30061), .ZN(I39767) );
INV_X32 U_g30308 ( .A(I39767), .ZN(g30308) );
INV_X32 U_I39770 ( .A(g30063), .ZN(I39770) );
INV_X32 U_g30309 ( .A(I39770), .ZN(g30309) );
INV_X32 U_I39773 ( .A(g30064), .ZN(I39773) );
INV_X32 U_g30310 ( .A(I39773), .ZN(g30310) );
INV_X32 U_I39776 ( .A(g30066), .ZN(I39776) );
INV_X32 U_g30311 ( .A(I39776), .ZN(g30311) );
INV_X32 U_I39779 ( .A(g30053), .ZN(I39779) );
INV_X32 U_g30312 ( .A(I39779), .ZN(g30312) );
INV_X32 U_I39782 ( .A(g30054), .ZN(I39782) );
INV_X32 U_g30313 ( .A(I39782), .ZN(g30313) );
INV_X32 U_I39785 ( .A(g30124), .ZN(I39785) );
INV_X32 U_g30314 ( .A(I39785), .ZN(g30314) );
INV_X32 U_I39788 ( .A(g30125), .ZN(I39788) );
INV_X32 U_g30315 ( .A(I39788), .ZN(g30315) );
INV_X32 U_I39791 ( .A(g30126), .ZN(I39791) );
INV_X32 U_g30316 ( .A(I39791), .ZN(g30316) );
INV_X32 U_I39794 ( .A(g30130), .ZN(I39794) );
INV_X32 U_g30317 ( .A(I39794), .ZN(g30317) );
INV_X32 U_I39797 ( .A(g30307), .ZN(I39797) );
INV_X32 U_g30318 ( .A(I39797), .ZN(g30318) );
INV_X32 U_I39800 ( .A(g30309), .ZN(I39800) );
INV_X32 U_g30319 ( .A(I39800), .ZN(g30319) );
INV_X32 U_I39803 ( .A(g30308), .ZN(I39803) );
INV_X32 U_g30320 ( .A(I39803), .ZN(g30320) );
INV_X32 U_I39806 ( .A(g30310), .ZN(I39806) );
INV_X32 U_g30321 ( .A(I39806), .ZN(g30321) );
INV_X32 U_I39809 ( .A(g30311), .ZN(I39809) );
INV_X32 U_g30322 ( .A(I39809), .ZN(g30322) );
INV_X32 U_I39812 ( .A(g30312), .ZN(I39812) );
INV_X32 U_g30323 ( .A(I39812), .ZN(g30323) );
INV_X32 U_I39815 ( .A(g30313), .ZN(I39815) );
INV_X32 U_g30324 ( .A(I39815), .ZN(g30324) );
INV_X32 U_I39818 ( .A(g30215), .ZN(I39818) );
INV_X32 U_g30325 ( .A(I39818), .ZN(g30325) );
INV_X32 U_I39821 ( .A(g30267), .ZN(I39821) );
INV_X32 U_g30326 ( .A(I39821), .ZN(g30326) );
INV_X32 U_I39825 ( .A(g30268), .ZN(I39825) );
INV_X32 U_g30328 ( .A(I39825), .ZN(g30328) );
INV_X32 U_I39828 ( .A(g30269), .ZN(I39828) );
INV_X32 U_g30329 ( .A(I39828), .ZN(g30329) );
INV_X32 U_I39832 ( .A(g30270), .ZN(I39832) );
INV_X32 U_g30331 ( .A(I39832), .ZN(g30331) );
INV_X32 U_I39835 ( .A(g30271), .ZN(I39835) );
INV_X32 U_g30332 ( .A(I39835), .ZN(g30332) );
INV_X32 U_I39840 ( .A(g30272), .ZN(I39840) );
INV_X32 U_g30335 ( .A(I39840), .ZN(g30335) );
INV_X32 U_I39843 ( .A(g30273), .ZN(I39843) );
INV_X32 U_g30336 ( .A(I39843), .ZN(g30336) );
INV_X32 U_I39848 ( .A(g30274), .ZN(I39848) );
INV_X32 U_g30339 ( .A(I39848), .ZN(g30339) );
INV_X32 U_I39853 ( .A(g30275), .ZN(I39853) );
INV_X32 U_g30342 ( .A(I39853), .ZN(g30342) );
INV_X32 U_I39856 ( .A(g30276), .ZN(I39856) );
INV_X32 U_g30343 ( .A(I39856), .ZN(g30343) );
INV_X32 U_I39859 ( .A(g30277), .ZN(I39859) );
INV_X32 U_g30344 ( .A(I39859), .ZN(g30344) );
INV_X32 U_I39863 ( .A(g30278), .ZN(I39863) );
INV_X32 U_g30346 ( .A(I39863), .ZN(g30346) );
INV_X32 U_I39866 ( .A(g30279), .ZN(I39866) );
INV_X32 U_g30347 ( .A(I39866), .ZN(g30347) );
INV_X32 U_I39870 ( .A(g30280), .ZN(I39870) );
INV_X32 U_g30349 ( .A(I39870), .ZN(g30349) );
INV_X32 U_I39873 ( .A(g30281), .ZN(I39873) );
INV_X32 U_g30350 ( .A(I39873), .ZN(g30350) );
INV_X32 U_I39878 ( .A(g30282), .ZN(I39878) );
INV_X32 U_g30353 ( .A(I39878), .ZN(g30353) );
INV_X32 U_I39881 ( .A(g30283), .ZN(I39881) );
INV_X32 U_g30354 ( .A(I39881), .ZN(g30354) );
INV_X32 U_I39886 ( .A(g30284), .ZN(I39886) );
INV_X32 U_g30357 ( .A(I39886), .ZN(g30357) );
INV_X32 U_I39889 ( .A(g30285), .ZN(I39889) );
INV_X32 U_g30358 ( .A(I39889), .ZN(g30358) );
INV_X32 U_I39892 ( .A(g30286), .ZN(I39892) );
INV_X32 U_g30359 ( .A(I39892), .ZN(g30359) );
INV_X32 U_I39895 ( .A(g30287), .ZN(I39895) );
INV_X32 U_g30360 ( .A(I39895), .ZN(g30360) );
INV_X32 U_I39899 ( .A(g30288), .ZN(I39899) );
INV_X32 U_g30362 ( .A(I39899), .ZN(g30362) );
INV_X32 U_I39902 ( .A(g30289), .ZN(I39902) );
INV_X32 U_g30363 ( .A(I39902), .ZN(g30363) );
INV_X32 U_I39906 ( .A(g30290), .ZN(I39906) );
INV_X32 U_g30365 ( .A(I39906), .ZN(g30365) );
INV_X32 U_I39909 ( .A(g30291), .ZN(I39909) );
INV_X32 U_g30366 ( .A(I39909), .ZN(g30366) );
INV_X32 U_I39913 ( .A(g30292), .ZN(I39913) );
INV_X32 U_g30368 ( .A(I39913), .ZN(g30368) );
INV_X32 U_I39916 ( .A(g30293), .ZN(I39916) );
INV_X32 U_g30369 ( .A(I39916), .ZN(g30369) );
INV_X32 U_I39919 ( .A(g30294), .ZN(I39919) );
INV_X32 U_g30370 ( .A(I39919), .ZN(g30370) );
INV_X32 U_I39922 ( .A(g30295), .ZN(I39922) );
INV_X32 U_g30371 ( .A(I39922), .ZN(g30371) );
INV_X32 U_I39926 ( .A(g30296), .ZN(I39926) );
INV_X32 U_g30373 ( .A(I39926), .ZN(g30373) );
INV_X32 U_I39930 ( .A(g30297), .ZN(I39930) );
INV_X32 U_g30375 ( .A(I39930), .ZN(g30375) );
INV_X32 U_I39933 ( .A(g30298), .ZN(I39933) );
INV_X32 U_g30376 ( .A(I39933), .ZN(g30376) );
INV_X32 U_I39936 ( .A(g30299), .ZN(I39936) );
INV_X32 U_g30377 ( .A(I39936), .ZN(g30377) );
INV_X32 U_I39939 ( .A(g30300), .ZN(I39939) );
INV_X32 U_g30378 ( .A(I39939), .ZN(g30378) );
INV_X32 U_I39942 ( .A(g30301), .ZN(I39942) );
INV_X32 U_g30379 ( .A(I39942), .ZN(g30379) );
INV_X32 U_I39945 ( .A(g30302), .ZN(I39945) );
INV_X32 U_g30380 ( .A(I39945), .ZN(g30380) );
INV_X32 U_I39948 ( .A(g30303), .ZN(I39948) );
INV_X32 U_g30381 ( .A(I39948), .ZN(g30381) );
INV_X32 U_I39951 ( .A(g30304), .ZN(I39951) );
INV_X32 U_g30382 ( .A(I39951), .ZN(g30382) );
INV_X32 U_g30383 ( .A(g30306), .ZN(g30383) );
INV_X32 U_I39976 ( .A(g30245), .ZN(I39976) );
INV_X32 U_g30408 ( .A(I39976), .ZN(g30408) );
INV_X32 U_I39982 ( .A(g30305), .ZN(I39982) );
INV_X32 U_g30412 ( .A(I39982), .ZN(g30412) );
INV_X32 U_I39985 ( .A(g30246), .ZN(I39985) );
INV_X32 U_g30435 ( .A(I39985), .ZN(g30435) );
INV_X32 U_I39991 ( .A(g30247), .ZN(I39991) );
INV_X32 U_g30439 ( .A(I39991), .ZN(g30439) );
INV_X32 U_I39997 ( .A(g30248), .ZN(I39997) );
INV_X32 U_g30443 ( .A(I39997), .ZN(g30443) );
INV_X32 U_I40002 ( .A(g30249), .ZN(I40002) );
INV_X32 U_g30446 ( .A(I40002), .ZN(g30446) );
INV_X32 U_I40008 ( .A(g30250), .ZN(I40008) );
INV_X32 U_g30450 ( .A(I40008), .ZN(g30450) );
INV_X32 U_I40016 ( .A(g30251), .ZN(I40016) );
INV_X32 U_g30456 ( .A(I40016), .ZN(g30456) );
INV_X32 U_I40021 ( .A(g30252), .ZN(I40021) );
INV_X32 U_g30459 ( .A(I40021), .ZN(g30459) );
INV_X32 U_I40027 ( .A(g30253), .ZN(I40027) );
INV_X32 U_g30463 ( .A(I40027), .ZN(g30463) );
INV_X32 U_I40032 ( .A(g30254), .ZN(I40032) );
INV_X32 U_g30466 ( .A(I40032), .ZN(g30466) );
INV_X32 U_I40039 ( .A(g30255), .ZN(I40039) );
INV_X32 U_g30471 ( .A(I40039), .ZN(g30471) );
INV_X32 U_I40044 ( .A(g30256), .ZN(I40044) );
INV_X32 U_g30474 ( .A(I40044), .ZN(g30474) );
INV_X32 U_I40051 ( .A(g30257), .ZN(I40051) );
INV_X32 U_g30479 ( .A(I40051), .ZN(g30479) );
INV_X32 U_I40054 ( .A(g30258), .ZN(I40054) );
INV_X32 U_g30480 ( .A(I40054), .ZN(g30480) );
INV_X32 U_I40059 ( .A(g30259), .ZN(I40059) );
INV_X32 U_g30483 ( .A(I40059), .ZN(g30483) );
INV_X32 U_I40066 ( .A(g30260), .ZN(I40066) );
INV_X32 U_g30488 ( .A(I40066), .ZN(g30488) );
INV_X32 U_I40071 ( .A(g30261), .ZN(I40071) );
INV_X32 U_g30491 ( .A(I40071), .ZN(g30491) );
INV_X32 U_I40075 ( .A(g30262), .ZN(I40075) );
INV_X32 U_g30493 ( .A(I40075), .ZN(g30493) );
INV_X32 U_I40078 ( .A(g30263), .ZN(I40078) );
INV_X32 U_g30494 ( .A(I40078), .ZN(g30494) );
INV_X32 U_I40083 ( .A(g30264), .ZN(I40083) );
INV_X32 U_g30497 ( .A(I40083), .ZN(g30497) );
INV_X32 U_I40086 ( .A(g30265), .ZN(I40086) );
INV_X32 U_g30498 ( .A(I40086), .ZN(g30498) );
INV_X32 U_I40091 ( .A(g30266), .ZN(I40091) );
INV_X32 U_g30501 ( .A(I40091), .ZN(g30501) );
INV_X32 U_I40098 ( .A(g30491), .ZN(I40098) );
INV_X32 U_g30506 ( .A(I40098), .ZN(g30506) );
INV_X32 U_I40101 ( .A(g30326), .ZN(I40101) );
INV_X32 U_g30507 ( .A(I40101), .ZN(g30507) );
INV_X32 U_I40104 ( .A(g30342), .ZN(I40104) );
INV_X32 U_g30508 ( .A(I40104), .ZN(g30508) );
INV_X32 U_I40107 ( .A(g30343), .ZN(I40107) );
INV_X32 U_g30509 ( .A(I40107), .ZN(g30509) );
INV_X32 U_I40110 ( .A(g30357), .ZN(I40110) );
INV_X32 U_g30510 ( .A(I40110), .ZN(g30510) );
INV_X32 U_I40113 ( .A(g30368), .ZN(I40113) );
INV_X32 U_g30511 ( .A(I40113), .ZN(g30511) );
INV_X32 U_I40116 ( .A(g30408), .ZN(I40116) );
INV_X32 U_g30512 ( .A(I40116), .ZN(g30512) );
INV_X32 U_I40119 ( .A(g30435), .ZN(I40119) );
INV_X32 U_g30513 ( .A(I40119), .ZN(g30513) );
INV_X32 U_I40122 ( .A(g30443), .ZN(I40122) );
INV_X32 U_g30514 ( .A(I40122), .ZN(g30514) );
INV_X32 U_I40125 ( .A(g30466), .ZN(I40125) );
INV_X32 U_g30515 ( .A(I40125), .ZN(g30515) );
INV_X32 U_I40128 ( .A(g30479), .ZN(I40128) );
INV_X32 U_g30516 ( .A(I40128), .ZN(g30516) );
INV_X32 U_I40131 ( .A(g30493), .ZN(I40131) );
INV_X32 U_g30517 ( .A(I40131), .ZN(g30517) );
INV_X32 U_I40134 ( .A(g30480), .ZN(I40134) );
INV_X32 U_g30518 ( .A(I40134), .ZN(g30518) );
INV_X32 U_I40137 ( .A(g30494), .ZN(I40137) );
INV_X32 U_g30519 ( .A(I40137), .ZN(g30519) );
INV_X32 U_I40140 ( .A(g30328), .ZN(I40140) );
INV_X32 U_g30520 ( .A(I40140), .ZN(g30520) );
INV_X32 U_I40143 ( .A(g30329), .ZN(I40143) );
INV_X32 U_g30521 ( .A(I40143), .ZN(g30521) );
INV_X32 U_I40146 ( .A(g30344), .ZN(I40146) );
INV_X32 U_g30522 ( .A(I40146), .ZN(g30522) );
INV_X32 U_I40149 ( .A(g30358), .ZN(I40149) );
INV_X32 U_g30523 ( .A(I40149), .ZN(g30523) );
INV_X32 U_I40152 ( .A(g30359), .ZN(I40152) );
INV_X32 U_g30524 ( .A(I40152), .ZN(g30524) );
INV_X32 U_I40155 ( .A(g30369), .ZN(I40155) );
INV_X32 U_g30525 ( .A(I40155), .ZN(g30525) );
INV_X32 U_I40158 ( .A(g30376), .ZN(I40158) );
INV_X32 U_g30526 ( .A(I40158), .ZN(g30526) );
INV_X32 U_I40161 ( .A(g30439), .ZN(I40161) );
INV_X32 U_g30527 ( .A(I40161), .ZN(g30527) );
INV_X32 U_I40164 ( .A(g30446), .ZN(I40164) );
INV_X32 U_g30528 ( .A(I40164), .ZN(g30528) );
INV_X32 U_I40167 ( .A(g30456), .ZN(I40167) );
INV_X32 U_g30529 ( .A(I40167), .ZN(g30529) );
INV_X32 U_I40170 ( .A(g30483), .ZN(I40170) );
INV_X32 U_g30530 ( .A(I40170), .ZN(g30530) );
INV_X32 U_I40173 ( .A(g30497), .ZN(I40173) );
INV_X32 U_g30531 ( .A(I40173), .ZN(g30531) );
INV_X32 U_I40176 ( .A(g30331), .ZN(I40176) );
INV_X32 U_g30532 ( .A(I40176), .ZN(g30532) );
INV_X32 U_I40179 ( .A(g30498), .ZN(I40179) );
INV_X32 U_g30533 ( .A(I40179), .ZN(g30533) );
INV_X32 U_I40182 ( .A(g30332), .ZN(I40182) );
INV_X32 U_g30534 ( .A(I40182), .ZN(g30534) );
INV_X32 U_I40185 ( .A(g30346), .ZN(I40185) );
INV_X32 U_g30535 ( .A(I40185), .ZN(g30535) );
INV_X32 U_I40188 ( .A(g30347), .ZN(I40188) );
INV_X32 U_g30536 ( .A(I40188), .ZN(g30536) );
INV_X32 U_I40191 ( .A(g30360), .ZN(I40191) );
INV_X32 U_g30537 ( .A(I40191), .ZN(g30537) );
INV_X32 U_I40194 ( .A(g30370), .ZN(I40194) );
INV_X32 U_g30538 ( .A(I40194), .ZN(g30538) );
INV_X32 U_I40197 ( .A(g30371), .ZN(I40197) );
INV_X32 U_g30539 ( .A(I40197), .ZN(g30539) );
INV_X32 U_I40200 ( .A(g30377), .ZN(I40200) );
INV_X32 U_g30540 ( .A(I40200), .ZN(g30540) );
INV_X32 U_I40203 ( .A(g30380), .ZN(I40203) );
INV_X32 U_g30541 ( .A(I40203), .ZN(g30541) );
INV_X32 U_I40206 ( .A(g30450), .ZN(I40206) );
INV_X32 U_g30542 ( .A(I40206), .ZN(g30542) );
INV_X32 U_I40209 ( .A(g30459), .ZN(I40209) );
INV_X32 U_g30543 ( .A(I40209), .ZN(g30543) );
INV_X32 U_I40212 ( .A(g30471), .ZN(I40212) );
INV_X32 U_g30544 ( .A(I40212), .ZN(g30544) );
INV_X32 U_I40215 ( .A(g30501), .ZN(I40215) );
INV_X32 U_g30545 ( .A(I40215), .ZN(g30545) );
INV_X32 U_I40218 ( .A(g30335), .ZN(I40218) );
INV_X32 U_g30546 ( .A(I40218), .ZN(g30546) );
INV_X32 U_I40221 ( .A(g30349), .ZN(I40221) );
INV_X32 U_g30547 ( .A(I40221), .ZN(g30547) );
INV_X32 U_I40224 ( .A(g30336), .ZN(I40224) );
INV_X32 U_g30548 ( .A(I40224), .ZN(g30548) );
INV_X32 U_I40227 ( .A(g30350), .ZN(I40227) );
INV_X32 U_g30549 ( .A(I40227), .ZN(g30549) );
INV_X32 U_I40230 ( .A(g30362), .ZN(I40230) );
INV_X32 U_g30550 ( .A(I40230), .ZN(g30550) );
INV_X32 U_I40233 ( .A(g30363), .ZN(I40233) );
INV_X32 U_g30551 ( .A(I40233), .ZN(g30551) );
INV_X32 U_I40236 ( .A(g30373), .ZN(I40236) );
INV_X32 U_g30552 ( .A(I40236), .ZN(g30552) );
INV_X32 U_I40239 ( .A(g30378), .ZN(I40239) );
INV_X32 U_g30553 ( .A(I40239), .ZN(g30553) );
INV_X32 U_I40242 ( .A(g30379), .ZN(I40242) );
INV_X32 U_g30554 ( .A(I40242), .ZN(g30554) );
INV_X32 U_I40245 ( .A(g30381), .ZN(I40245) );
INV_X32 U_g30555 ( .A(I40245), .ZN(g30555) );
INV_X32 U_I40248 ( .A(g30382), .ZN(I40248) );
INV_X32 U_g30556 ( .A(I40248), .ZN(g30556) );
INV_X32 U_I40251 ( .A(g30463), .ZN(I40251) );
INV_X32 U_g30557 ( .A(I40251), .ZN(g30557) );
INV_X32 U_I40254 ( .A(g30474), .ZN(I40254) );
INV_X32 U_g30558 ( .A(I40254), .ZN(g30558) );
INV_X32 U_I40257 ( .A(g30488), .ZN(I40257) );
INV_X32 U_g30559 ( .A(I40257), .ZN(g30559) );
INV_X32 U_I40260 ( .A(g30339), .ZN(I40260) );
INV_X32 U_g30560 ( .A(I40260), .ZN(g30560) );
INV_X32 U_I40263 ( .A(g30353), .ZN(I40263) );
INV_X32 U_g30561 ( .A(I40263), .ZN(g30561) );
INV_X32 U_I40266 ( .A(g30365), .ZN(I40266) );
INV_X32 U_g30562 ( .A(I40266), .ZN(g30562) );
INV_X32 U_I40269 ( .A(g30354), .ZN(I40269) );
INV_X32 U_g30563 ( .A(I40269), .ZN(g30563) );
INV_X32 U_I40272 ( .A(g30366), .ZN(I40272) );
INV_X32 U_g30564 ( .A(I40272), .ZN(g30564) );
INV_X32 U_I40275 ( .A(g30375), .ZN(I40275) );
INV_X32 U_g30565 ( .A(I40275), .ZN(g30565) );
INV_X32 U_g30567 ( .A(g30403), .ZN(g30567) );
INV_X32 U_g30568 ( .A(g30402), .ZN(g30568) );
INV_X32 U_g30569 ( .A(g30406), .ZN(g30569) );
INV_X32 U_g30570 ( .A(g30404), .ZN(g30570) );
INV_X32 U_g30571 ( .A(g30401), .ZN(g30571) );
INV_X32 U_g30572 ( .A(g30399), .ZN(g30572) );
INV_X32 U_g30573 ( .A(g30405), .ZN(g30573) );
INV_X32 U_g30574 ( .A(g30400), .ZN(g30574) );
INV_X32 U_g30575 ( .A(g30412), .ZN(g30575) );
INV_X32 U_I40288 ( .A(g30455), .ZN(I40288) );
INV_X32 U_g30578 ( .A(I40288), .ZN(g30578) );
INV_X32 U_I40291 ( .A(g30468), .ZN(I40291) );
INV_X32 U_g30579 ( .A(I40291), .ZN(g30579) );
INV_X32 U_I40294 ( .A(g30470), .ZN(I40294) );
INV_X32 U_g30580 ( .A(I40294), .ZN(g30580) );
INV_X32 U_I40297 ( .A(g30482), .ZN(I40297) );
INV_X32 U_g30581 ( .A(I40297), .ZN(g30581) );
INV_X32 U_I40300 ( .A(g30485), .ZN(I40300) );
INV_X32 U_g30582 ( .A(I40300), .ZN(g30582) );
INV_X32 U_I40303 ( .A(g30487), .ZN(I40303) );
INV_X32 U_g30583 ( .A(I40303), .ZN(g30583) );
INV_X32 U_I40307 ( .A(g30500), .ZN(I40307) );
INV_X32 U_g30585 ( .A(I40307), .ZN(g30585) );
INV_X32 U_I40310 ( .A(g30503), .ZN(I40310) );
INV_X32 U_g30586 ( .A(I40310), .ZN(g30586) );
INV_X32 U_I40313 ( .A(g30505), .ZN(I40313) );
INV_X32 U_g30587 ( .A(I40313), .ZN(g30587) );
INV_X32 U_I40317 ( .A(g30338), .ZN(I40317) );
INV_X32 U_g30591 ( .A(I40317), .ZN(g30591) );
INV_X32 U_I40320 ( .A(g30341), .ZN(I40320) );
INV_X32 U_g30592 ( .A(I40320), .ZN(g30592) );
INV_X32 U_I40326 ( .A(g30356), .ZN(I40326) );
INV_X32 U_g30600 ( .A(I40326), .ZN(g30600) );
INV_X32 U_I40420 ( .A(g30578), .ZN(I40420) );
INV_X32 U_g30710 ( .A(I40420), .ZN(g30710) );
INV_X32 U_I40423 ( .A(g30579), .ZN(I40423) );
INV_X32 U_g30711 ( .A(I40423), .ZN(g30711) );
INV_X32 U_I40426 ( .A(g30581), .ZN(I40426) );
INV_X32 U_g30712 ( .A(I40426), .ZN(g30712) );
INV_X32 U_I40429 ( .A(g30580), .ZN(I40429) );
INV_X32 U_g30713 ( .A(I40429), .ZN(g30713) );
INV_X32 U_I40432 ( .A(g30582), .ZN(I40432) );
INV_X32 U_g30714 ( .A(I40432), .ZN(g30714) );
INV_X32 U_I40435 ( .A(g30585), .ZN(I40435) );
INV_X32 U_g30715 ( .A(I40435), .ZN(g30715) );
INV_X32 U_I40438 ( .A(g30583), .ZN(I40438) );
INV_X32 U_g30716 ( .A(I40438), .ZN(g30716) );
INV_X32 U_I40441 ( .A(g30586), .ZN(I40441) );
INV_X32 U_g30717 ( .A(I40441), .ZN(g30717) );
INV_X32 U_I40444 ( .A(g30591), .ZN(I40444) );
INV_X32 U_g30718 ( .A(I40444), .ZN(g30718) );
INV_X32 U_I40447 ( .A(g30587), .ZN(I40447) );
INV_X32 U_g30719 ( .A(I40447), .ZN(g30719) );
INV_X32 U_I40450 ( .A(g30592), .ZN(I40450) );
INV_X32 U_g30720 ( .A(I40450), .ZN(g30720) );
INV_X32 U_I40453 ( .A(g30600), .ZN(I40453) );
INV_X32 U_g30721 ( .A(I40453), .ZN(g30721) );
INV_X32 U_I40456 ( .A(g30668), .ZN(I40456) );
INV_X32 U_g30722 ( .A(I40456), .ZN(g30722) );
INV_X32 U_I40459 ( .A(g30669), .ZN(I40459) );
INV_X32 U_g30723 ( .A(I40459), .ZN(g30723) );
INV_X32 U_I40462 ( .A(g30670), .ZN(I40462) );
INV_X32 U_g30724 ( .A(I40462), .ZN(g30724) );
INV_X32 U_I40465 ( .A(g30671), .ZN(I40465) );
INV_X32 U_g30725 ( .A(I40465), .ZN(g30725) );
INV_X32 U_I40468 ( .A(g30672), .ZN(I40468) );
INV_X32 U_g30726 ( .A(I40468), .ZN(g30726) );
INV_X32 U_I40471 ( .A(g30673), .ZN(I40471) );
INV_X32 U_g30727 ( .A(I40471), .ZN(g30727) );
INV_X32 U_I40475 ( .A(g30674), .ZN(I40475) );
INV_X32 U_g30729 ( .A(I40475), .ZN(g30729) );
INV_X32 U_I40478 ( .A(g30675), .ZN(I40478) );
INV_X32 U_g30730 ( .A(I40478), .ZN(g30730) );
INV_X32 U_I40481 ( .A(g30676), .ZN(I40481) );
INV_X32 U_g30731 ( .A(I40481), .ZN(g30731) );
INV_X32 U_I40484 ( .A(g30677), .ZN(I40484) );
INV_X32 U_g30732 ( .A(I40484), .ZN(g30732) );
INV_X32 U_I40487 ( .A(g30678), .ZN(I40487) );
INV_X32 U_g30733 ( .A(I40487), .ZN(g30733) );
INV_X32 U_I40490 ( .A(g30679), .ZN(I40490) );
INV_X32 U_g30734 ( .A(I40490), .ZN(g30734) );
INV_X32 U_I40495 ( .A(g30680), .ZN(I40495) );
INV_X32 U_g30737 ( .A(I40495), .ZN(g30737) );
INV_X32 U_I40498 ( .A(g30681), .ZN(I40498) );
INV_X32 U_g30738 ( .A(I40498), .ZN(g30738) );
INV_X32 U_I40501 ( .A(g30682), .ZN(I40501) );
INV_X32 U_g30739 ( .A(I40501), .ZN(g30739) );
INV_X32 U_I40504 ( .A(g30683), .ZN(I40504) );
INV_X32 U_g30740 ( .A(I40504), .ZN(g30740) );
INV_X32 U_I40507 ( .A(g30684), .ZN(I40507) );
INV_X32 U_g30741 ( .A(I40507), .ZN(g30741) );
INV_X32 U_I40510 ( .A(g30686), .ZN(I40510) );
INV_X32 U_g30742 ( .A(I40510), .ZN(g30742) );
INV_X32 U_I40515 ( .A(g30687), .ZN(I40515) );
INV_X32 U_g30745 ( .A(I40515), .ZN(g30745) );
INV_X32 U_I40518 ( .A(g30688), .ZN(I40518) );
INV_X32 U_g30746 ( .A(I40518), .ZN(g30746) );
INV_X32 U_I40521 ( .A(g30689), .ZN(I40521) );
INV_X32 U_g30747 ( .A(I40521), .ZN(g30747) );
INV_X32 U_I40524 ( .A(g30690), .ZN(I40524) );
INV_X32 U_g30748 ( .A(I40524), .ZN(g30748) );
INV_X32 U_I40527 ( .A(g30691), .ZN(I40527) );
INV_X32 U_g30749 ( .A(I40527), .ZN(g30749) );
INV_X32 U_I40531 ( .A(g30692), .ZN(I40531) );
INV_X32 U_g30751 ( .A(I40531), .ZN(g30751) );
INV_X32 U_I40534 ( .A(g30693), .ZN(I40534) );
INV_X32 U_g30752 ( .A(I40534), .ZN(g30752) );
INV_X32 U_I40537 ( .A(g30694), .ZN(I40537) );
INV_X32 U_g30753 ( .A(I40537), .ZN(g30753) );
INV_X32 U_I40542 ( .A(g30695), .ZN(I40542) );
INV_X32 U_g30756 ( .A(I40542), .ZN(g30756) );
INV_X32 U_g30765 ( .A(g30685), .ZN(g30765) );
INV_X32 U_I40555 ( .A(g30699), .ZN(I40555) );
INV_X32 U_g30767 ( .A(I40555), .ZN(g30767) );
INV_X32 U_I40565 ( .A(g30700), .ZN(I40565) );
INV_X32 U_g30769 ( .A(I40565), .ZN(g30769) );
INV_X32 U_I40568 ( .A(g30701), .ZN(I40568) );
INV_X32 U_g30770 ( .A(I40568), .ZN(g30770) );
INV_X32 U_I40578 ( .A(g30702), .ZN(I40578) );
INV_X32 U_g30772 ( .A(I40578), .ZN(g30772) );
INV_X32 U_I40581 ( .A(g30703), .ZN(I40581) );
INV_X32 U_g30773 ( .A(I40581), .ZN(g30773) );
INV_X32 U_I40584 ( .A(g30704), .ZN(I40584) );
INV_X32 U_g30774 ( .A(I40584), .ZN(g30774) );
INV_X32 U_I40594 ( .A(g30705), .ZN(I40594) );
INV_X32 U_g30776 ( .A(I40594), .ZN(g30776) );
INV_X32 U_I40597 ( .A(g30706), .ZN(I40597) );
INV_X32 U_g30777 ( .A(I40597), .ZN(g30777) );
INV_X32 U_I40600 ( .A(g30707), .ZN(I40600) );
INV_X32 U_g30778 ( .A(I40600), .ZN(g30778) );
INV_X32 U_I40611 ( .A(g30708), .ZN(I40611) );
INV_X32 U_g30781 ( .A(I40611), .ZN(g30781) );
INV_X32 U_I40614 ( .A(g30709), .ZN(I40614) );
INV_X32 U_g30782 ( .A(I40614), .ZN(g30782) );
INV_X32 U_I40618 ( .A(g30566), .ZN(I40618) );
INV_X32 U_g30784 ( .A(I40618), .ZN(g30784) );
INV_X32 U_I40634 ( .A(g30571), .ZN(I40634) );
INV_X32 U_g30792 ( .A(I40634), .ZN(g30792) );
INV_X32 U_I40637 ( .A(g30570), .ZN(I40637) );
INV_X32 U_g30793 ( .A(I40637), .ZN(g30793) );
INV_X32 U_I40640 ( .A(g30569), .ZN(I40640) );
INV_X32 U_g30794 ( .A(I40640), .ZN(g30794) );
INV_X32 U_I40643 ( .A(g30568), .ZN(I40643) );
INV_X32 U_g30795 ( .A(I40643), .ZN(g30795) );
INV_X32 U_I40647 ( .A(g30567), .ZN(I40647) );
INV_X32 U_g30797 ( .A(I40647), .ZN(g30797) );
INV_X32 U_I40651 ( .A(g30574), .ZN(I40651) );
INV_X32 U_g30799 ( .A(I40651), .ZN(g30799) );
INV_X32 U_I40654 ( .A(g30573), .ZN(I40654) );
INV_X32 U_g30800 ( .A(I40654), .ZN(g30800) );
INV_X32 U_I40658 ( .A(g30572), .ZN(I40658) );
INV_X32 U_g30802 ( .A(I40658), .ZN(g30802) );
INV_X32 U_I40661 ( .A(g30635), .ZN(I40661) );
INV_X32 U_g30803 ( .A(I40661), .ZN(g30803) );
INV_X32 U_I40664 ( .A(g30636), .ZN(I40664) );
INV_X32 U_g30804 ( .A(I40664), .ZN(g30804) );
INV_X32 U_I40667 ( .A(g30637), .ZN(I40667) );
INV_X32 U_g30805 ( .A(I40667), .ZN(g30805) );
INV_X32 U_I40670 ( .A(g30638), .ZN(I40670) );
INV_X32 U_g30806 ( .A(I40670), .ZN(g30806) );
INV_X32 U_I40673 ( .A(g30639), .ZN(I40673) );
INV_X32 U_g30807 ( .A(I40673), .ZN(g30807) );
INV_X32 U_I40676 ( .A(g30640), .ZN(I40676) );
INV_X32 U_g30808 ( .A(I40676), .ZN(g30808) );
INV_X32 U_I40679 ( .A(g30641), .ZN(I40679) );
INV_X32 U_g30809 ( .A(I40679), .ZN(g30809) );
INV_X32 U_I40682 ( .A(g30642), .ZN(I40682) );
INV_X32 U_g30810 ( .A(I40682), .ZN(g30810) );
INV_X32 U_I40685 ( .A(g30643), .ZN(I40685) );
INV_X32 U_g30811 ( .A(I40685), .ZN(g30811) );
INV_X32 U_I40688 ( .A(g30644), .ZN(I40688) );
INV_X32 U_g30812 ( .A(I40688), .ZN(g30812) );
INV_X32 U_I40691 ( .A(g30645), .ZN(I40691) );
INV_X32 U_g30813 ( .A(I40691), .ZN(g30813) );
INV_X32 U_I40694 ( .A(g30646), .ZN(I40694) );
INV_X32 U_g30814 ( .A(I40694), .ZN(g30814) );
INV_X32 U_I40697 ( .A(g30647), .ZN(I40697) );
INV_X32 U_g30815 ( .A(I40697), .ZN(g30815) );
INV_X32 U_I40700 ( .A(g30648), .ZN(I40700) );
INV_X32 U_g30816 ( .A(I40700), .ZN(g30816) );
INV_X32 U_I40703 ( .A(g30649), .ZN(I40703) );
INV_X32 U_g30817 ( .A(I40703), .ZN(g30817) );
INV_X32 U_I40706 ( .A(g30650), .ZN(I40706) );
INV_X32 U_g30818 ( .A(I40706), .ZN(g30818) );
INV_X32 U_I40709 ( .A(g30651), .ZN(I40709) );
INV_X32 U_g30819 ( .A(I40709), .ZN(g30819) );
INV_X32 U_I40712 ( .A(g30652), .ZN(I40712) );
INV_X32 U_g30820 ( .A(I40712), .ZN(g30820) );
INV_X32 U_I40715 ( .A(g30653), .ZN(I40715) );
INV_X32 U_g30821 ( .A(I40715), .ZN(g30821) );
INV_X32 U_I40718 ( .A(g30654), .ZN(I40718) );
INV_X32 U_g30822 ( .A(I40718), .ZN(g30822) );
INV_X32 U_I40721 ( .A(g30655), .ZN(I40721) );
INV_X32 U_g30823 ( .A(I40721), .ZN(g30823) );
INV_X32 U_I40724 ( .A(g30656), .ZN(I40724) );
INV_X32 U_g30824 ( .A(I40724), .ZN(g30824) );
INV_X32 U_I40727 ( .A(g30657), .ZN(I40727) );
INV_X32 U_g30825 ( .A(I40727), .ZN(g30825) );
INV_X32 U_I40730 ( .A(g30658), .ZN(I40730) );
INV_X32 U_g30826 ( .A(I40730), .ZN(g30826) );
INV_X32 U_I40733 ( .A(g30659), .ZN(I40733) );
INV_X32 U_g30827 ( .A(I40733), .ZN(g30827) );
INV_X32 U_I40736 ( .A(g30660), .ZN(I40736) );
INV_X32 U_g30828 ( .A(I40736), .ZN(g30828) );
INV_X32 U_I40739 ( .A(g30661), .ZN(I40739) );
INV_X32 U_g30829 ( .A(I40739), .ZN(g30829) );
INV_X32 U_I40742 ( .A(g30662), .ZN(I40742) );
INV_X32 U_g30830 ( .A(I40742), .ZN(g30830) );
INV_X32 U_I40745 ( .A(g30663), .ZN(I40745) );
INV_X32 U_g30831 ( .A(I40745), .ZN(g30831) );
INV_X32 U_I40748 ( .A(g30664), .ZN(I40748) );
INV_X32 U_g30832 ( .A(I40748), .ZN(g30832) );
INV_X32 U_I40751 ( .A(g30665), .ZN(I40751) );
INV_X32 U_g30833 ( .A(I40751), .ZN(g30833) );
INV_X32 U_I40754 ( .A(g30666), .ZN(I40754) );
INV_X32 U_g30834 ( .A(I40754), .ZN(g30834) );
INV_X32 U_I40757 ( .A(g30667), .ZN(I40757) );
INV_X32 U_g30835 ( .A(I40757), .ZN(g30835) );
INV_X32 U_I40760 ( .A(g30722), .ZN(I40760) );
INV_X32 U_g30836 ( .A(I40760), .ZN(g30836) );
INV_X32 U_I40763 ( .A(g30729), .ZN(I40763) );
INV_X32 U_g30837 ( .A(I40763), .ZN(g30837) );
INV_X32 U_I40766 ( .A(g30737), .ZN(I40766) );
INV_X32 U_g30838 ( .A(I40766), .ZN(g30838) );
INV_X32 U_I40769 ( .A(g30803), .ZN(I40769) );
INV_X32 U_g30839 ( .A(I40769), .ZN(g30839) );
INV_X32 U_I40772 ( .A(g30804), .ZN(I40772) );
INV_X32 U_g30840 ( .A(I40772), .ZN(g30840) );
INV_X32 U_I40775 ( .A(g30807), .ZN(I40775) );
INV_X32 U_g30841 ( .A(I40775), .ZN(g30841) );
INV_X32 U_I40778 ( .A(g30805), .ZN(I40778) );
INV_X32 U_g30842 ( .A(I40778), .ZN(g30842) );
INV_X32 U_I40781 ( .A(g30808), .ZN(I40781) );
INV_X32 U_g30843 ( .A(I40781), .ZN(g30843) );
INV_X32 U_I40784 ( .A(g30813), .ZN(I40784) );
INV_X32 U_g30844 ( .A(I40784), .ZN(g30844) );
INV_X32 U_I40787 ( .A(g30809), .ZN(I40787) );
INV_X32 U_g30845 ( .A(I40787), .ZN(g30845) );
INV_X32 U_I40790 ( .A(g30814), .ZN(I40790) );
INV_X32 U_g30846 ( .A(I40790), .ZN(g30846) );
INV_X32 U_I40793 ( .A(g30821), .ZN(I40793) );
INV_X32 U_g30847 ( .A(I40793), .ZN(g30847) );
INV_X32 U_I40796 ( .A(g30829), .ZN(I40796) );
INV_X32 U_g30848 ( .A(I40796), .ZN(g30848) );
INV_X32 U_I40799 ( .A(g30723), .ZN(I40799) );
INV_X32 U_g30849 ( .A(I40799), .ZN(g30849) );
INV_X32 U_I40802 ( .A(g30730), .ZN(I40802) );
INV_X32 U_g30850 ( .A(I40802), .ZN(g30850) );
INV_X32 U_I40805 ( .A(g30767), .ZN(I40805) );
INV_X32 U_g30851 ( .A(I40805), .ZN(g30851) );
INV_X32 U_I40808 ( .A(g30769), .ZN(I40808) );
INV_X32 U_g30852 ( .A(I40808), .ZN(g30852) );
INV_X32 U_I40811 ( .A(g30772), .ZN(I40811) );
INV_X32 U_g30853 ( .A(I40811), .ZN(g30853) );
INV_X32 U_I40814 ( .A(g30731), .ZN(I40814) );
INV_X32 U_g30854 ( .A(I40814), .ZN(g30854) );
INV_X32 U_I40817 ( .A(g30738), .ZN(I40817) );
INV_X32 U_g30855 ( .A(I40817), .ZN(g30855) );
INV_X32 U_I40820 ( .A(g30745), .ZN(I40820) );
INV_X32 U_g30856 ( .A(I40820), .ZN(g30856) );
INV_X32 U_I40823 ( .A(g30806), .ZN(I40823) );
INV_X32 U_g30857 ( .A(I40823), .ZN(g30857) );
INV_X32 U_I40826 ( .A(g30810), .ZN(I40826) );
INV_X32 U_g30858 ( .A(I40826), .ZN(g30858) );
INV_X32 U_I40829 ( .A(g30815), .ZN(I40829) );
INV_X32 U_g30859 ( .A(I40829), .ZN(g30859) );
INV_X32 U_I40832 ( .A(g30811), .ZN(I40832) );
INV_X32 U_g30860 ( .A(I40832), .ZN(g30860) );
INV_X32 U_I40835 ( .A(g30816), .ZN(I40835) );
INV_X32 U_g30861 ( .A(I40835), .ZN(g30861) );
INV_X32 U_I40838 ( .A(g30822), .ZN(I40838) );
INV_X32 U_g30862 ( .A(I40838), .ZN(g30862) );
INV_X32 U_I40841 ( .A(g30817), .ZN(I40841) );
INV_X32 U_g30863 ( .A(I40841), .ZN(g30863) );
INV_X32 U_I40844 ( .A(g30823), .ZN(I40844) );
INV_X32 U_g30864 ( .A(I40844), .ZN(g30864) );
INV_X32 U_I40847 ( .A(g30830), .ZN(I40847) );
INV_X32 U_g30865 ( .A(I40847), .ZN(g30865) );
INV_X32 U_I40850 ( .A(g30724), .ZN(I40850) );
INV_X32 U_g30866 ( .A(I40850), .ZN(g30866) );
INV_X32 U_I40853 ( .A(g30732), .ZN(I40853) );
INV_X32 U_g30867 ( .A(I40853), .ZN(g30867) );
INV_X32 U_I40856 ( .A(g30739), .ZN(I40856) );
INV_X32 U_g30868 ( .A(I40856), .ZN(g30868) );
INV_X32 U_I40859 ( .A(g30770), .ZN(I40859) );
INV_X32 U_g30869 ( .A(I40859), .ZN(g30869) );
INV_X32 U_I40862 ( .A(g30773), .ZN(I40862) );
INV_X32 U_g30870 ( .A(I40862), .ZN(g30870) );
INV_X32 U_I40865 ( .A(g30776), .ZN(I40865) );
INV_X32 U_g30871 ( .A(I40865), .ZN(g30871) );
INV_X32 U_I40868 ( .A(g30740), .ZN(I40868) );
INV_X32 U_g30872 ( .A(I40868), .ZN(g30872) );
INV_X32 U_I40871 ( .A(g30746), .ZN(I40871) );
INV_X32 U_g30873 ( .A(I40871), .ZN(g30873) );
INV_X32 U_I40874 ( .A(g30751), .ZN(I40874) );
INV_X32 U_g30874 ( .A(I40874), .ZN(g30874) );
INV_X32 U_I40877 ( .A(g30812), .ZN(I40877) );
INV_X32 U_g30875 ( .A(I40877), .ZN(g30875) );
INV_X32 U_I40880 ( .A(g30818), .ZN(I40880) );
INV_X32 U_g30876 ( .A(I40880), .ZN(g30876) );
INV_X32 U_I40883 ( .A(g30824), .ZN(I40883) );
INV_X32 U_g30877 ( .A(I40883), .ZN(g30877) );
INV_X32 U_I40886 ( .A(g30819), .ZN(I40886) );
INV_X32 U_g30878 ( .A(I40886), .ZN(g30878) );
INV_X32 U_I40889 ( .A(g30825), .ZN(I40889) );
INV_X32 U_g30879 ( .A(I40889), .ZN(g30879) );
INV_X32 U_I40892 ( .A(g30831), .ZN(I40892) );
INV_X32 U_g30880 ( .A(I40892), .ZN(g30880) );
INV_X32 U_I40895 ( .A(g30826), .ZN(I40895) );
INV_X32 U_g30881 ( .A(I40895), .ZN(g30881) );
INV_X32 U_I40898 ( .A(g30832), .ZN(I40898) );
INV_X32 U_g30882 ( .A(I40898), .ZN(g30882) );
INV_X32 U_I40901 ( .A(g30725), .ZN(I40901) );
INV_X32 U_g30883 ( .A(I40901), .ZN(g30883) );
INV_X32 U_I40904 ( .A(g30733), .ZN(I40904) );
INV_X32 U_g30884 ( .A(I40904), .ZN(g30884) );
INV_X32 U_I40907 ( .A(g30741), .ZN(I40907) );
INV_X32 U_g30885 ( .A(I40907), .ZN(g30885) );
INV_X32 U_I40910 ( .A(g30747), .ZN(I40910) );
INV_X32 U_g30886 ( .A(I40910), .ZN(g30886) );
INV_X32 U_I40913 ( .A(g30774), .ZN(I40913) );
INV_X32 U_g30887 ( .A(I40913), .ZN(g30887) );
INV_X32 U_I40916 ( .A(g30777), .ZN(I40916) );
INV_X32 U_g30888 ( .A(I40916), .ZN(g30888) );
INV_X32 U_I40919 ( .A(g30781), .ZN(I40919) );
INV_X32 U_g30889 ( .A(I40919), .ZN(g30889) );
INV_X32 U_I40922 ( .A(g30748), .ZN(I40922) );
INV_X32 U_g30890 ( .A(I40922), .ZN(g30890) );
INV_X32 U_I40925 ( .A(g30752), .ZN(I40925) );
INV_X32 U_g30891 ( .A(I40925), .ZN(g30891) );
INV_X32 U_I40928 ( .A(g30756), .ZN(I40928) );
INV_X32 U_g30892 ( .A(I40928), .ZN(g30892) );
INV_X32 U_I40931 ( .A(g30820), .ZN(I40931) );
INV_X32 U_g30893 ( .A(I40931), .ZN(g30893) );
INV_X32 U_I40934 ( .A(g30827), .ZN(I40934) );
INV_X32 U_g30894 ( .A(I40934), .ZN(g30894) );
INV_X32 U_I40937 ( .A(g30833), .ZN(I40937) );
INV_X32 U_g30895 ( .A(I40937), .ZN(g30895) );
INV_X32 U_I40940 ( .A(g30828), .ZN(I40940) );
INV_X32 U_g30896 ( .A(I40940), .ZN(g30896) );
INV_X32 U_I40943 ( .A(g30834), .ZN(I40943) );
INV_X32 U_g30897 ( .A(I40943), .ZN(g30897) );
INV_X32 U_I40946 ( .A(g30726), .ZN(I40946) );
INV_X32 U_g30898 ( .A(I40946), .ZN(g30898) );
INV_X32 U_I40949 ( .A(g30835), .ZN(I40949) );
INV_X32 U_g30899 ( .A(I40949), .ZN(g30899) );
INV_X32 U_I40952 ( .A(g30727), .ZN(I40952) );
INV_X32 U_g30900 ( .A(I40952), .ZN(g30900) );
INV_X32 U_I40955 ( .A(g30734), .ZN(I40955) );
INV_X32 U_g30901 ( .A(I40955), .ZN(g30901) );
INV_X32 U_I40958 ( .A(g30742), .ZN(I40958) );
INV_X32 U_g30902 ( .A(I40958), .ZN(g30902) );
INV_X32 U_I40961 ( .A(g30749), .ZN(I40961) );
INV_X32 U_g30903 ( .A(I40961), .ZN(g30903) );
INV_X32 U_I40964 ( .A(g30753), .ZN(I40964) );
INV_X32 U_g30904 ( .A(I40964), .ZN(g30904) );
INV_X32 U_I40967 ( .A(g30778), .ZN(I40967) );
INV_X32 U_g30905 ( .A(I40967), .ZN(g30905) );
INV_X32 U_I40970 ( .A(g30782), .ZN(I40970) );
INV_X32 U_g30906 ( .A(I40970), .ZN(g30906) );
INV_X32 U_I40973 ( .A(g30784), .ZN(I40973) );
INV_X32 U_g30907 ( .A(I40973), .ZN(g30907) );
INV_X32 U_I40976 ( .A(g30799), .ZN(I40976) );
INV_X32 U_g30908 ( .A(I40976), .ZN(g30908) );
INV_X32 U_I40979 ( .A(g30800), .ZN(I40979) );
INV_X32 U_g30909 ( .A(I40979), .ZN(g30909) );
INV_X32 U_I40982 ( .A(g30802), .ZN(I40982) );
INV_X32 U_g30910 ( .A(I40982), .ZN(g30910) );
INV_X32 U_I40985 ( .A(g30792), .ZN(I40985) );
INV_X32 U_g30911 ( .A(I40985), .ZN(g30911) );
INV_X32 U_I40988 ( .A(g30793), .ZN(I40988) );
INV_X32 U_g30912 ( .A(I40988), .ZN(g30912) );
INV_X32 U_I40991 ( .A(g30794), .ZN(I40991) );
INV_X32 U_g30913 ( .A(I40991), .ZN(g30913) );
INV_X32 U_I40994 ( .A(g30795), .ZN(I40994) );
INV_X32 U_g30914 ( .A(I40994), .ZN(g30914) );
INV_X32 U_I40997 ( .A(g30797), .ZN(I40997) );
INV_X32 U_g30915 ( .A(I40997), .ZN(g30915) );
INV_X32 U_I41024 ( .A(g30765), .ZN(I41024) );
INV_X32 U_g30928 ( .A(I41024), .ZN(g30928) );
INV_X32 U_I41035 ( .A(g30796), .ZN(I41035) );
INV_X32 U_g30937 ( .A(I41035), .ZN(g30937) );
INV_X32 U_I41038 ( .A(g30798), .ZN(I41038) );
INV_X32 U_g30938 ( .A(I41038), .ZN(g30938) );
INV_X32 U_I41041 ( .A(g30801), .ZN(I41041) );
INV_X32 U_g30939 ( .A(I41041), .ZN(g30939) );
INV_X32 U_I41044 ( .A(g30928), .ZN(I41044) );
INV_X32 U_g30940 ( .A(I41044), .ZN(g30940) );
INV_X32 U_I41047 ( .A(g30937), .ZN(I41047) );
INV_X32 U_g30941 ( .A(I41047), .ZN(g30941) );
INV_X32 U_I41050 ( .A(g30938), .ZN(I41050) );
INV_X32 U_g30942 ( .A(I41050), .ZN(g30942) );
INV_X32 U_I41053 ( .A(g30939), .ZN(I41053) );
INV_X32 U_g30943 ( .A(I41053), .ZN(g30943) );
INV_X32 U_g30962 ( .A(g30958), .ZN(g30962) );
INV_X32 U_g30963 ( .A(g30957), .ZN(g30963) );
INV_X32 U_g30964 ( .A(g30961), .ZN(g30964) );
INV_X32 U_g30965 ( .A(g30959), .ZN(g30965) );
INV_X32 U_g30966 ( .A(g30956), .ZN(g30966) );
INV_X32 U_g30967 ( .A(g30954), .ZN(g30967) );
INV_X32 U_g30968 ( .A(g30960), .ZN(g30968) );
INV_X32 U_g30969 ( .A(g30955), .ZN(g30969) );
INV_X32 U_g30971 ( .A(g30970), .ZN(g30971) );
INV_X32 U_I41090 ( .A(g30965), .ZN(I41090) );
INV_X32 U_g30972 ( .A(I41090), .ZN(g30972) );
INV_X32 U_I41093 ( .A(g30964), .ZN(I41093) );
INV_X32 U_g30973 ( .A(I41093), .ZN(g30973) );
INV_X32 U_I41096 ( .A(g30963), .ZN(I41096) );
INV_X32 U_g30974 ( .A(I41096), .ZN(g30974) );
INV_X32 U_I41099 ( .A(g30962), .ZN(I41099) );
INV_X32 U_g30975 ( .A(I41099), .ZN(g30975) );
INV_X32 U_I41102 ( .A(g30969), .ZN(I41102) );
INV_X32 U_g30976 ( .A(I41102), .ZN(g30976) );
INV_X32 U_I41105 ( .A(g30968), .ZN(I41105) );
INV_X32 U_g30977 ( .A(I41105), .ZN(g30977) );
INV_X32 U_I41108 ( .A(g30967), .ZN(I41108) );
INV_X32 U_g30978 ( .A(I41108), .ZN(g30978) );
INV_X32 U_I41111 ( .A(g30966), .ZN(I41111) );
INV_X32 U_g30979 ( .A(I41111), .ZN(g30979) );
INV_X32 U_I41114 ( .A(g30976), .ZN(I41114) );
INV_X32 U_g30980 ( .A(I41114), .ZN(g30980) );
INV_X32 U_I41117 ( .A(g30977), .ZN(I41117) );
INV_X32 U_g30981 ( .A(I41117), .ZN(g30981) );
INV_X32 U_I41120 ( .A(g30978), .ZN(I41120) );
INV_X32 U_g30982 ( .A(I41120), .ZN(g30982) );
INV_X32 U_I41123 ( .A(g30979), .ZN(I41123) );
INV_X32 U_g30983 ( .A(I41123), .ZN(g30983) );
INV_X32 U_I41126 ( .A(g30972), .ZN(I41126) );
INV_X32 U_g30984 ( .A(I41126), .ZN(g30984) );
INV_X32 U_I41129 ( .A(g30973), .ZN(I41129) );
INV_X32 U_g30985 ( .A(I41129), .ZN(g30985) );
INV_X32 U_I41132 ( .A(g30974), .ZN(I41132) );
INV_X32 U_g30986 ( .A(I41132), .ZN(g30986) );
INV_X32 U_I41135 ( .A(g30975), .ZN(I41135) );
INV_X32 U_g30987 ( .A(I41135), .ZN(g30987) );
INV_X32 U_I41138 ( .A(g30971), .ZN(I41138) );
INV_X32 U_g30988 ( .A(I41138), .ZN(g30988) );
INV_X32 U_I41141 ( .A(g30988), .ZN(I41141) );
INV_X32 U_g30989 ( .A(I41141), .ZN(g30989) );
AND2_X4 U_g5630 ( .A1(g325), .A2(g349), .ZN(g5630) );
AND2_X4 U_g5649 ( .A1(g331), .A2(g351), .ZN(g5649) );
AND2_X4 U_g5650 ( .A1(g325), .A2(g364), .ZN(g5650) );
AND2_X4 U_g5658 ( .A1(g1012), .A2(g1036), .ZN(g5658) );
AND2_X4 U_g5676 ( .A1(g337), .A2(g353), .ZN(g5676) );
AND2_X4 U_g5677 ( .A1(g331), .A2(g366), .ZN(g5677) );
AND2_X4 U_g5678 ( .A1(g325), .A2(g379), .ZN(g5678) );
AND2_X4 U_g5687 ( .A1(g1018), .A2(g1038), .ZN(g5687) );
AND2_X4 U_g5688 ( .A1(g1012), .A2(g1051), .ZN(g5688) );
AND2_X4 U_g5696 ( .A1(g1706), .A2(g1730), .ZN(g5696) );
AND2_X4 U_g5709 ( .A1(g337), .A2(g368), .ZN(g5709) );
AND2_X4 U_g5710 ( .A1(g331), .A2(g381), .ZN(g5710) );
AND2_X4 U_g5711 ( .A1(g325), .A2(g394), .ZN(g5711) );
AND2_X4 U_g5728 ( .A1(g1024), .A2(g1040), .ZN(g5728) );
AND2_X4 U_g5729 ( .A1(g1018), .A2(g1053), .ZN(g5729) );
AND2_X4 U_g5730 ( .A1(g1012), .A2(g1066), .ZN(g5730) );
AND2_X4 U_g5739 ( .A1(g1712), .A2(g1732), .ZN(g5739) );
AND2_X4 U_g5740 ( .A1(g1706), .A2(g1745), .ZN(g5740) );
AND2_X4 U_g5748 ( .A1(g2400), .A2(g2424), .ZN(g5748) );
AND2_X4 U_g5757 ( .A1(g337), .A2(g383), .ZN(g5757) );
AND2_X4 U_g5758 ( .A1(g331), .A2(g396), .ZN(g5758) );
AND2_X4 U_g5767 ( .A1(g1024), .A2(g1055), .ZN(g5767) );
AND2_X4 U_g5768 ( .A1(g1018), .A2(g1068), .ZN(g5768) );
AND2_X4 U_g5769 ( .A1(g1012), .A2(g1081), .ZN(g5769) );
AND2_X4 U_g5786 ( .A1(g1718), .A2(g1734), .ZN(g5786) );
AND2_X4 U_g5787 ( .A1(g1712), .A2(g1747), .ZN(g5787) );
AND2_X4 U_g5788 ( .A1(g1706), .A2(g1760), .ZN(g5788) );
AND2_X4 U_g5797 ( .A1(g2406), .A2(g2426), .ZN(g5797) );
AND2_X4 U_g5798 ( .A1(g2400), .A2(g2439), .ZN(g5798) );
AND2_X4 U_g5807 ( .A1(g337), .A2(g324), .ZN(g5807) );
AND2_X4 U_g5816 ( .A1(g1024), .A2(g1070), .ZN(g5816) );
AND2_X4 U_g5817 ( .A1(g1018), .A2(g1083), .ZN(g5817) );
AND2_X4 U_g5826 ( .A1(g1718), .A2(g1749), .ZN(g5826) );
AND2_X4 U_g5827 ( .A1(g1712), .A2(g1762), .ZN(g5827) );
AND2_X4 U_g5828 ( .A1(g1706), .A2(g1775), .ZN(g5828) );
AND2_X4 U_g5845 ( .A1(g2412), .A2(g2428), .ZN(g5845) );
AND2_X4 U_g5846 ( .A1(g2406), .A2(g2441), .ZN(g5846) );
AND2_X4 U_g5847 ( .A1(g2400), .A2(g2454), .ZN(g5847) );
AND2_X4 U_g5863 ( .A1(g1024), .A2(g1011), .ZN(g5863) );
AND2_X4 U_g5872 ( .A1(g1718), .A2(g1764), .ZN(g5872) );
AND2_X4 U_g5873 ( .A1(g1712), .A2(g1777), .ZN(g5873) );
AND2_X4 U_g5882 ( .A1(g2412), .A2(g2443), .ZN(g5882) );
AND2_X4 U_g5883 ( .A1(g2406), .A2(g2456), .ZN(g5883) );
AND2_X4 U_g5884 ( .A1(g2400), .A2(g2469), .ZN(g5884) );
AND2_X4 U_g5910 ( .A1(g1718), .A2(g1705), .ZN(g5910) );
AND2_X4 U_g5919 ( .A1(g2412), .A2(g2458), .ZN(g5919) );
AND2_X4 U_g5920 ( .A1(g2406), .A2(g2471), .ZN(g5920) );
AND2_X4 U_g5949 ( .A1(g2412), .A2(g2399), .ZN(g5949) );
AND2_X4 U_g8327 ( .A1(g3254), .A2(g219), .ZN(g8327) );
AND2_X4 U_g8328 ( .A1(g6314), .A2(g225), .ZN(g8328) );
AND2_X4 U_g8329 ( .A1(g6232), .A2(g231), .ZN(g8329) );
AND2_X4 U_g8339 ( .A1(g6519), .A2(g903), .ZN(g8339) );
AND2_X4 U_g8340 ( .A1(g6369), .A2(g909), .ZN(g8340) );
AND2_X4 U_g8350 ( .A1(g6574), .A2(g1594), .ZN(g8350) );
AND2_X4 U_g8385 ( .A1(g3254), .A2(g228), .ZN(g8385) );
AND2_X4 U_g8386 ( .A1(g6314), .A2(g234), .ZN(g8386) );
AND2_X4 U_g8387 ( .A1(g6232), .A2(g240), .ZN(g8387) );
AND2_X4 U_g8394 ( .A1(g3410), .A2(g906), .ZN(g8394) );
AND2_X4 U_g8395 ( .A1(g6519), .A2(g912), .ZN(g8395) );
AND2_X4 U_g8396 ( .A1(g6369), .A2(g918), .ZN(g8396) );
AND2_X4 U_g8406 ( .A1(g6783), .A2(g1597), .ZN(g8406) );
AND2_X4 U_g8407 ( .A1(g6574), .A2(g1603), .ZN(g8407) );
AND2_X4 U_g8417 ( .A1(g6838), .A2(g2288), .ZN(g8417) );
AND2_X4 U_g8431 ( .A1(g3254), .A2(g237), .ZN(g8431) );
AND2_X4 U_g8432 ( .A1(g6314), .A2(g243), .ZN(g8432) );
AND2_X4 U_g8433 ( .A1(g6232), .A2(g249), .ZN(g8433) );
AND2_X4 U_g8437 ( .A1(g3410), .A2(g915), .ZN(g8437) );
AND2_X4 U_g8438 ( .A1(g6519), .A2(g921), .ZN(g8438) );
AND2_X4 U_g8439 ( .A1(g6369), .A2(g927), .ZN(g8439) );
AND2_X4 U_g8446 ( .A1(g3566), .A2(g1600), .ZN(g8446) );
AND2_X4 U_g8447 ( .A1(g6783), .A2(g1606), .ZN(g8447) );
AND2_X4 U_g8448 ( .A1(g6574), .A2(g1612), .ZN(g8448) );
AND2_X4 U_g8458 ( .A1(g7085), .A2(g2291), .ZN(g8458) );
AND2_X4 U_g8459 ( .A1(g6838), .A2(g2297), .ZN(g8459) );
AND2_X4 U_g8463 ( .A1(g3254), .A2(g246), .ZN(g8463) );
AND2_X4 U_g8464 ( .A1(g6314), .A2(g252), .ZN(g8464) );
AND2_X4 U_g8465 ( .A1(g6232), .A2(g258), .ZN(g8465) );
AND2_X4 U_g8466 ( .A1(g3410), .A2(g924), .ZN(g8466) );
AND2_X4 U_g8467 ( .A1(g6519), .A2(g930), .ZN(g8467) );
AND2_X4 U_g8468 ( .A1(g6369), .A2(g936), .ZN(g8468) );
AND2_X4 U_g8472 ( .A1(g3566), .A2(g1609), .ZN(g8472) );
AND2_X4 U_g8473 ( .A1(g6783), .A2(g1615), .ZN(g8473) );
AND2_X4 U_g8474 ( .A1(g6574), .A2(g1621), .ZN(g8474) );
AND2_X4 U_g8481 ( .A1(g3722), .A2(g2294), .ZN(g8481) );
AND2_X4 U_g8482 ( .A1(g7085), .A2(g2300), .ZN(g8482) );
AND2_X4 U_g8483 ( .A1(g6838), .A2(g2306), .ZN(g8483) );
AND2_X4 U_g8484 ( .A1(g6232), .A2(g186), .ZN(g8484) );
AND2_X4 U_g8485 ( .A1(g3254), .A2(g255), .ZN(g8485) );
AND2_X4 U_g8486 ( .A1(g6314), .A2(g261), .ZN(g8486) );
AND2_X4 U_g8487 ( .A1(g6232), .A2(g267), .ZN(g8487) );
AND2_X4 U_g8488 ( .A1(g3410), .A2(g933), .ZN(g8488) );
AND2_X4 U_g8489 ( .A1(g6519), .A2(g939), .ZN(g8489) );
AND2_X4 U_g8490 ( .A1(g6369), .A2(g945), .ZN(g8490) );
AND2_X4 U_g8491 ( .A1(g3566), .A2(g1618), .ZN(g8491) );
AND2_X4 U_g8492 ( .A1(g6783), .A2(g1624), .ZN(g8492) );
AND2_X4 U_g8493 ( .A1(g6574), .A2(g1630), .ZN(g8493) );
AND2_X4 U_g8497 ( .A1(g3722), .A2(g2303), .ZN(g8497) );
AND2_X4 U_g8498 ( .A1(g7085), .A2(g2309), .ZN(g8498) );
AND2_X4 U_g8499 ( .A1(g6838), .A2(g2315), .ZN(g8499) );
AND2_X4 U_g8500 ( .A1(g6314), .A2(g189), .ZN(g8500) );
AND2_X4 U_g8501 ( .A1(g6232), .A2(g195), .ZN(g8501) );
AND2_X4 U_g8502 ( .A1(g3254), .A2(g264), .ZN(g8502) );
AND2_X4 U_g8503 ( .A1(g6314), .A2(g270), .ZN(g8503) );
AND2_X4 U_g8504 ( .A1(g6369), .A2(g873), .ZN(g8504) );
AND2_X4 U_g8505 ( .A1(g3410), .A2(g942), .ZN(g8505) );
AND2_X4 U_g8506 ( .A1(g6519), .A2(g948), .ZN(g8506) );
AND2_X4 U_g8507 ( .A1(g6369), .A2(g954), .ZN(g8507) );
AND2_X4 U_g8508 ( .A1(g3566), .A2(g1627), .ZN(g8508) );
AND2_X4 U_g8509 ( .A1(g6783), .A2(g1633), .ZN(g8509) );
AND2_X4 U_g8510 ( .A1(g6574), .A2(g1639), .ZN(g8510) );
AND2_X4 U_g8511 ( .A1(g3722), .A2(g2312), .ZN(g8511) );
AND2_X4 U_g8512 ( .A1(g7085), .A2(g2318), .ZN(g8512) );
AND2_X4 U_g8513 ( .A1(g6838), .A2(g2324), .ZN(g8513) );
AND2_X4 U_g8515 ( .A1(g3254), .A2(g192), .ZN(g8515) );
AND2_X4 U_g8516 ( .A1(g6314), .A2(g198), .ZN(g8516) );
AND2_X4 U_g8517 ( .A1(g6232), .A2(g204), .ZN(g8517) );
AND2_X4 U_g8518 ( .A1(g3254), .A2(g273), .ZN(g8518) );
AND2_X4 U_g8519 ( .A1(g6519), .A2(g876), .ZN(g8519) );
AND2_X4 U_g8520 ( .A1(g6369), .A2(g882), .ZN(g8520) );
AND2_X4 U_g8521 ( .A1(g3410), .A2(g951), .ZN(g8521) );
AND2_X4 U_g8522 ( .A1(g6519), .A2(g957), .ZN(g8522) );
AND2_X4 U_g8523 ( .A1(g6574), .A2(g1567), .ZN(g8523) );
AND2_X4 U_g8524 ( .A1(g3566), .A2(g1636), .ZN(g8524) );
AND2_X4 U_g8525 ( .A1(g6783), .A2(g1642), .ZN(g8525) );
AND2_X4 U_g8526 ( .A1(g6574), .A2(g1648), .ZN(g8526) );
AND2_X4 U_g8527 ( .A1(g3722), .A2(g2321), .ZN(g8527) );
AND2_X4 U_g8528 ( .A1(g7085), .A2(g2327), .ZN(g8528) );
AND2_X4 U_g8529 ( .A1(g6838), .A2(g2333), .ZN(g8529) );
AND2_X4 U_g8531 ( .A1(g3254), .A2(g201), .ZN(g8531) );
AND2_X4 U_g8532 ( .A1(g6314), .A2(g207), .ZN(g8532) );
AND2_X4 U_g8534 ( .A1(g3410), .A2(g879), .ZN(g8534) );
AND2_X4 U_g8535 ( .A1(g6519), .A2(g885), .ZN(g8535) );
AND2_X4 U_g8536 ( .A1(g6369), .A2(g891), .ZN(g8536) );
AND2_X4 U_g8537 ( .A1(g3410), .A2(g960), .ZN(g8537) );
AND2_X4 U_g8538 ( .A1(g6783), .A2(g1570), .ZN(g8538) );
AND2_X4 U_g8539 ( .A1(g6574), .A2(g1576), .ZN(g8539) );
AND2_X4 U_g8540 ( .A1(g3566), .A2(g1645), .ZN(g8540) );
AND2_X4 U_g8541 ( .A1(g6783), .A2(g1651), .ZN(g8541) );
AND2_X4 U_g8542 ( .A1(g6838), .A2(g2261), .ZN(g8542) );
AND2_X4 U_g8543 ( .A1(g3722), .A2(g2330), .ZN(g8543) );
AND2_X4 U_g8544 ( .A1(g7085), .A2(g2336), .ZN(g8544) );
AND2_X4 U_g8545 ( .A1(g6838), .A2(g2342), .ZN(g8545) );
AND2_X4 U_g8546 ( .A1(g3254), .A2(g210), .ZN(g8546) );
AND2_X4 U_g8548 ( .A1(g3410), .A2(g888), .ZN(g8548) );
AND2_X4 U_g8549 ( .A1(g6519), .A2(g894), .ZN(g8549) );
AND2_X4 U_g8551 ( .A1(g3566), .A2(g1573), .ZN(g8551) );
AND2_X4 U_g8552 ( .A1(g6783), .A2(g1579), .ZN(g8552) );
AND2_X4 U_g8553 ( .A1(g6574), .A2(g1585), .ZN(g8553) );
AND2_X4 U_g8554 ( .A1(g3566), .A2(g1654), .ZN(g8554) );
AND2_X4 U_g8555 ( .A1(g7085), .A2(g2264), .ZN(g8555) );
AND2_X4 U_g8556 ( .A1(g6838), .A2(g2270), .ZN(g8556) );
AND2_X4 U_g8557 ( .A1(g3722), .A2(g2339), .ZN(g8557) );
AND2_X4 U_g8558 ( .A1(g7085), .A2(g2345), .ZN(g8558) );
AND2_X4 U_g8559 ( .A1(g3410), .A2(g897), .ZN(g8559) );
AND2_X4 U_g8561 ( .A1(g3566), .A2(g1582), .ZN(g8561) );
AND2_X4 U_g8562 ( .A1(g6783), .A2(g1588), .ZN(g8562) );
AND2_X4 U_g8564 ( .A1(g3722), .A2(g2267), .ZN(g8564) );
AND2_X4 U_g8565 ( .A1(g7085), .A2(g2273), .ZN(g8565) );
AND2_X4 U_g8566 ( .A1(g6838), .A2(g2279), .ZN(g8566) );
AND2_X4 U_g8567 ( .A1(g3722), .A2(g2348), .ZN(g8567) );
AND2_X4 U_g8570 ( .A1(g3566), .A2(g1591), .ZN(g8570) );
AND2_X4 U_g8572 ( .A1(g3722), .A2(g2276), .ZN(g8572) );
AND2_X4 U_g8573 ( .A1(g7085), .A2(g2282), .ZN(g8573) );
AND2_X4 U_g8576 ( .A1(g3722), .A2(g2285), .ZN(g8576) );
AND2_X4 U_g8601 ( .A1(g6643), .A2(g7153), .ZN(g8601) );
AND2_X4 U_g8612 ( .A1(g3338), .A2(g6908), .ZN(g8612) );
AND2_X4 U_g8613 ( .A1(g6945), .A2(g7349), .ZN(g8613) );
AND2_X4 U_g8621 ( .A1(g6486), .A2(g6672), .ZN(g8621) );
AND2_X4 U_g8625 ( .A1(g3494), .A2(g7158), .ZN(g8625) );
AND2_X4 U_g8626 ( .A1(g7195), .A2(g7479), .ZN(g8626) );
AND2_X4 U_g8631 ( .A1(g6751), .A2(g6974), .ZN(g8631) );
AND2_X4 U_g8635 ( .A1(g3650), .A2(g7354), .ZN(g8635) );
AND2_X4 U_g8636 ( .A1(g7391), .A2(g7535), .ZN(g8636) );
AND2_X4 U_g8650 ( .A1(g7053), .A2(g7224), .ZN(g8650) );
AND2_X4 U_g8654 ( .A1(g3806), .A2(g7484), .ZN(g8654) );
AND2_X4 U_g8666 ( .A1(g7303), .A2(g7420), .ZN(g8666) );
AND2_X4 U_g8676 ( .A1(g6643), .A2(g7838), .ZN(g8676) );
AND2_X4 U_g8687 ( .A1(g3338), .A2(g7827), .ZN(g8687) );
AND2_X4 U_g8688 ( .A1(g6945), .A2(g7858), .ZN(g8688) );
AND2_X4 U_g8703 ( .A1(g6486), .A2(g7819), .ZN(g8703) );
AND2_X4 U_g8704 ( .A1(g6643), .A2(g7996), .ZN(g8704) );
AND2_X4 U_g8705 ( .A1(g3494), .A2(g7842), .ZN(g8705) );
AND2_X4 U_g8706 ( .A1(g7195), .A2(g7888), .ZN(g8706) );
AND2_X4 U_g8717 ( .A1(g3338), .A2(g7953), .ZN(g8717) );
AND2_X4 U_g8722 ( .A1(g6751), .A2(g7830), .ZN(g8722) );
AND2_X4 U_g8723 ( .A1(g6945), .A2(g8071), .ZN(g8723) );
AND2_X4 U_g8724 ( .A1(g3650), .A2(g7862), .ZN(g8724) );
AND2_X4 U_g8725 ( .A1(g7391), .A2(g7912), .ZN(g8725) );
AND2_X4 U_g8751 ( .A1(g6486), .A2(g7906), .ZN(g8751) );
AND2_X4 U_g8755 ( .A1(g3494), .A2(g8004), .ZN(g8755) );
AND2_X4 U_g8760 ( .A1(g7053), .A2(g7845), .ZN(g8760) );
AND2_X4 U_g8761 ( .A1(g7195), .A2(g8156), .ZN(g8761) );
AND2_X4 U_g8762 ( .A1(g3806), .A2(g7892), .ZN(g8762) );
AND2_X4 U_g8774 ( .A1(g6751), .A2(g7958), .ZN(g8774) );
AND2_X4 U_g8778 ( .A1(g3650), .A2(g8079), .ZN(g8778) );
AND2_X4 U_g8783 ( .A1(g7303), .A2(g7865), .ZN(g8783) );
AND2_X4 U_g8784 ( .A1(g7391), .A2(g8242), .ZN(g8784) );
AND2_X4 U_g8797 ( .A1(g7053), .A2(g8009), .ZN(g8797) );
AND2_X4 U_g8801 ( .A1(g3806), .A2(g8164), .ZN(g8801) );
AND2_X4 U_g8816 ( .A1(g7303), .A2(g8084), .ZN(g8816) );
AND2_X4 U_g8841 ( .A1(g6486), .A2(g490), .ZN(g8841) );
AND2_X4 U_g8842 ( .A1(g6512), .A2(g5508), .ZN(g8842) );
AND2_X4 U_g8861 ( .A1(g6643), .A2(g493), .ZN(g8861) );
AND2_X4 U_g8868 ( .A1(g6751), .A2(g1177), .ZN(g8868) );
AND2_X4 U_g8869 ( .A1(g6776), .A2(g5552), .ZN(g8869) );
AND2_X4 U_g8892 ( .A1(g3338), .A2(g496), .ZN(g8892) );
AND2_X4 U_g8899 ( .A1(g6945), .A2(g1180), .ZN(g8899) );
AND2_X4 U_g8906 ( .A1(g7053), .A2(g1871), .ZN(g8906) );
AND2_X4 U_g8907 ( .A1(g7078), .A2(g5598), .ZN(g8907) );
AND2_X4 U_g8932 ( .A1(g3494), .A2(g1183), .ZN(g8932) );
AND2_X4 U_g8939 ( .A1(g7195), .A2(g1874), .ZN(g8939) );
AND2_X4 U_g8946 ( .A1(g7303), .A2(g2565), .ZN(g8946) );
AND2_X4 U_g8947 ( .A1(g7328), .A2(g5615), .ZN(g8947) );
AND2_X4 U_g8972 ( .A1(g3650), .A2(g1877), .ZN(g8972) );
AND2_X4 U_g8979 ( .A1(g7391), .A2(g2568), .ZN(g8979) );
AND2_X4 U_g9004 ( .A1(g3806), .A2(g2571), .ZN(g9004) );
AND2_X4 U_g9009 ( .A1(g6486), .A2(g565), .ZN(g9009) );
AND2_X4 U_g9026 ( .A1(g5438), .A2(g7610), .ZN(g9026) );
AND2_X4 U_g9033 ( .A1(g6643), .A2(g567), .ZN(g9033) );
AND2_X4 U_g9034 ( .A1(g6751), .A2(g1251), .ZN(g9034) );
AND2_X4 U_g9047 ( .A1(g6448), .A2(g7616), .ZN(g9047) );
AND2_X4 U_g9048 ( .A1(g3338), .A2(g489), .ZN(g9048) );
AND2_X4 U_g9049 ( .A1(g5473), .A2(g7619), .ZN(g9049) );
AND2_X4 U_g9056 ( .A1(g6945), .A2(g1253), .ZN(g9056) );
AND2_X4 U_g9057 ( .A1(g7053), .A2(g1945), .ZN(g9057) );
AND2_X4 U_g9061 ( .A1(g3306), .A2(g7623), .ZN(g9061) );
AND2_X4 U_g9062 ( .A1(g5438), .A2(g7626), .ZN(g9062) );
AND2_X4 U_g9063 ( .A1(g5438), .A2(g7629), .ZN(g9063) );
AND2_X4 U_g9064 ( .A1(g6713), .A2(g7632), .ZN(g9064) );
AND2_X4 U_g9065 ( .A1(g3494), .A2(g1176), .ZN(g9065) );
AND2_X4 U_g9066 ( .A1(g5512), .A2(g7635), .ZN(g9066) );
AND2_X4 U_g9073 ( .A1(g7195), .A2(g1947), .ZN(g9073) );
AND2_X4 U_g9074 ( .A1(g7303), .A2(g2639), .ZN(g9074) );
AND2_X4 U_g9075 ( .A1(g6448), .A2(g7643), .ZN(g9075) );
AND2_X4 U_g9076 ( .A1(g5438), .A2(g7646), .ZN(g9076) );
AND2_X4 U_g9077 ( .A1(g6448), .A2(g7649), .ZN(g9077) );
AND2_X4 U_g9078 ( .A1(g3462), .A2(g7652), .ZN(g9078) );
AND2_X4 U_g9079 ( .A1(g5473), .A2(g7655), .ZN(g9079) );
AND2_X4 U_g9080 ( .A1(g5473), .A2(g7658), .ZN(g9080) );
AND2_X4 U_g9081 ( .A1(g7015), .A2(g7661), .ZN(g9081) );
AND2_X4 U_g9082 ( .A1(g3650), .A2(g1870), .ZN(g9082) );
AND2_X4 U_g9083 ( .A1(g5556), .A2(g7664), .ZN(g9083) );
AND2_X4 U_g9090 ( .A1(g7391), .A2(g2641), .ZN(g9090) );
AND2_X4 U_g9091 ( .A1(g3306), .A2(g7670), .ZN(g9091) );
AND2_X4 U_g9092 ( .A1(g6448), .A2(g7673), .ZN(g9092) );
AND2_X4 U_g9093 ( .A1(g3306), .A2(g7676), .ZN(g9093) );
AND2_X4 U_g9094 ( .A1(g6713), .A2(g7679), .ZN(g9094) );
AND2_X4 U_g9095 ( .A1(g5473), .A2(g7682), .ZN(g9095) );
AND2_X4 U_g9096 ( .A1(g6713), .A2(g7685), .ZN(g9096) );
AND2_X4 U_g9097 ( .A1(g3618), .A2(g7688), .ZN(g9097) );
AND2_X4 U_g9098 ( .A1(g5512), .A2(g7691), .ZN(g9098) );
AND2_X4 U_g9099 ( .A1(g5512), .A2(g7694), .ZN(g9099) );
AND2_X4 U_g9100 ( .A1(g7265), .A2(g7697), .ZN(g9100) );
AND2_X4 U_g9101 ( .A1(g3806), .A2(g2564), .ZN(g9101) );
AND2_X4 U_g9102 ( .A1(g3306), .A2(g7703), .ZN(g9102) );
AND2_X4 U_g9103 ( .A1(g3462), .A2(g7706), .ZN(g9103) );
AND2_X4 U_g9104 ( .A1(g6713), .A2(g7709), .ZN(g9104) );
AND2_X4 U_g9105 ( .A1(g3462), .A2(g7712), .ZN(g9105) );
AND2_X4 U_g9106 ( .A1(g7015), .A2(g7715), .ZN(g9106) );
AND2_X4 U_g9107 ( .A1(g5512), .A2(g7718), .ZN(g9107) );
AND2_X4 U_g9108 ( .A1(g7015), .A2(g7721), .ZN(g9108) );
AND2_X4 U_g9109 ( .A1(g3774), .A2(g7724), .ZN(g9109) );
AND2_X4 U_g9110 ( .A1(g5556), .A2(g7727), .ZN(g9110) );
AND2_X4 U_g9111 ( .A1(g5556), .A2(g7730), .ZN(g9111) );
AND2_X4 U_g9112 ( .A1(g3462), .A2(g7733), .ZN(g9112) );
AND2_X4 U_g9113 ( .A1(g3618), .A2(g7736), .ZN(g9113) );
AND2_X4 U_g9114 ( .A1(g7015), .A2(g7739), .ZN(g9114) );
AND2_X4 U_g9115 ( .A1(g3618), .A2(g7742), .ZN(g9115) );
AND2_X4 U_g9116 ( .A1(g7265), .A2(g7745), .ZN(g9116) );
AND2_X4 U_g9117 ( .A1(g5556), .A2(g7748), .ZN(g9117) );
AND2_X4 U_g9118 ( .A1(g7265), .A2(g7751), .ZN(g9118) );
AND2_X4 U_g9119 ( .A1(g5438), .A2(g7754), .ZN(g9119) );
AND2_X4 U_g9120 ( .A1(g3618), .A2(g7757), .ZN(g9120) );
AND2_X4 U_g9121 ( .A1(g3774), .A2(g7760), .ZN(g9121) );
AND2_X4 U_g9122 ( .A1(g7265), .A2(g7763), .ZN(g9122) );
AND2_X4 U_g9123 ( .A1(g3774), .A2(g7766), .ZN(g9123) );
AND2_X4 U_g9124 ( .A1(g6448), .A2(g7769), .ZN(g9124) );
AND2_X4 U_g9125 ( .A1(g5473), .A2(g7776), .ZN(g9125) );
AND2_X4 U_g9126 ( .A1(g3774), .A2(g7779), .ZN(g9126) );
AND2_X4 U_g9127 ( .A1(g3306), .A2(g7782), .ZN(g9127) );
AND2_X4 U_g9131 ( .A1(g6713), .A2(g7785), .ZN(g9131) );
AND2_X4 U_g9132 ( .A1(g5512), .A2(g7792), .ZN(g9132) );
AND2_X4 U_g9133 ( .A1(g3462), .A2(g7796), .ZN(g9133) );
AND2_X4 U_g9137 ( .A1(g7015), .A2(g7799), .ZN(g9137) );
AND2_X4 U_g9138 ( .A1(g5556), .A2(g7806), .ZN(g9138) );
AND2_X4 U_g9139 ( .A1(g3618), .A2(g7809), .ZN(g9139) );
AND2_X4 U_g9143 ( .A1(g7265), .A2(g7812), .ZN(g9143) );
AND2_X4 U_g9145 ( .A1(g3774), .A2(g7823), .ZN(g9145) );
AND2_X4 U_g9241 ( .A1(g6232), .A2(g7950), .ZN(g9241) );
AND2_X4 U_g9301 ( .A1(g6314), .A2(g7990), .ZN(g9301) );
AND2_X4 U_g9302 ( .A1(g6232), .A2(g7993), .ZN(g9302) );
AND2_X4 U_g9319 ( .A1(g6369), .A2(g8001), .ZN(g9319) );
AND2_X4 U_g9364 ( .A1(g3254), .A2(g8053), .ZN(g9364) );
AND2_X4 U_g9365 ( .A1(g6314), .A2(g8056), .ZN(g9365) );
AND2_X4 U_g9366 ( .A1(g6232), .A2(g8059), .ZN(g9366) );
AND2_X4 U_g9367 ( .A1(g6232), .A2(g8062), .ZN(g9367) );
AND2_X4 U_g9382 ( .A1(g6519), .A2(g8065), .ZN(g9382) );
AND2_X4 U_g9383 ( .A1(g6369), .A2(g8068), .ZN(g9383) );
AND2_X4 U_g9400 ( .A1(g6574), .A2(g8076), .ZN(g9400) );
AND2_X4 U_g9438 ( .A1(g3254), .A2(g8123), .ZN(g9438) );
AND2_X4 U_g9439 ( .A1(g6314), .A2(g8126), .ZN(g9439) );
AND2_X4 U_g9440 ( .A1(g6232), .A2(g8129), .ZN(g9440) );
AND2_X4 U_g9441 ( .A1(g6314), .A2(g8132), .ZN(g9441) );
AND2_X4 U_g9442 ( .A1(g6232), .A2(g8135), .ZN(g9442) );
AND2_X4 U_g9461 ( .A1(g3410), .A2(g8138), .ZN(g9461) );
AND2_X4 U_g9462 ( .A1(g6519), .A2(g8141), .ZN(g9462) );
AND2_X4 U_g9463 ( .A1(g6369), .A2(g8144), .ZN(g9463) );
AND2_X4 U_g9464 ( .A1(g6369), .A2(g8147), .ZN(g9464) );
AND2_X4 U_g9479 ( .A1(g6783), .A2(g8150), .ZN(g9479) );
AND2_X4 U_g9480 ( .A1(g6574), .A2(g8153), .ZN(g9480) );
AND2_X4 U_g9497 ( .A1(g6838), .A2(g8161), .ZN(g9497) );
AND2_X4 U_g9518 ( .A1(g3254), .A2(g8191), .ZN(g9518) );
AND2_X4 U_g9519 ( .A1(g6314), .A2(g8194), .ZN(g9519) );
AND2_X4 U_g9520 ( .A1(g6232), .A2(g8197), .ZN(g9520) );
AND2_X4 U_g9521 ( .A1(g3254), .A2(g8200), .ZN(g9521) );
AND2_X4 U_g9522 ( .A1(g6314), .A2(g8203), .ZN(g9522) );
AND2_X4 U_g9523 ( .A1(g6232), .A2(g8206), .ZN(g9523) );
AND3_X4 U_g9534 ( .A1(g7772), .A2(g6135), .A3(g538), .ZN(g9534) );
AND2_X4 U_g9580 ( .A1(g3410), .A2(g8209), .ZN(g9580) );
AND2_X4 U_g9581 ( .A1(g6519), .A2(g8212), .ZN(g9581) );
AND2_X4 U_g9582 ( .A1(g6369), .A2(g8215), .ZN(g9582) );
AND2_X4 U_g9583 ( .A1(g6519), .A2(g8218), .ZN(g9583) );
AND2_X4 U_g9584 ( .A1(g6369), .A2(g8221), .ZN(g9584) );
AND2_X4 U_g9603 ( .A1(g3566), .A2(g8224), .ZN(g9603) );
AND2_X4 U_g9604 ( .A1(g6783), .A2(g8227), .ZN(g9604) );
AND2_X4 U_g9605 ( .A1(g6574), .A2(g8230), .ZN(g9605) );
AND2_X4 U_g9606 ( .A1(g6574), .A2(g8233), .ZN(g9606) );
AND2_X4 U_g9621 ( .A1(g7085), .A2(g8236), .ZN(g9621) );
AND2_X4 U_g9622 ( .A1(g6838), .A2(g8239), .ZN(g9622) );
AND2_X4 U_g9630 ( .A1(g3254), .A2(g3922), .ZN(g9630) );
AND2_X4 U_g9631 ( .A1(g6314), .A2(g3925), .ZN(g9631) );
AND2_X4 U_g9632 ( .A1(g6232), .A2(g3928), .ZN(g9632) );
AND2_X4 U_g9633 ( .A1(g3254), .A2(g3931), .ZN(g9633) );
AND2_X4 U_g9634 ( .A1(g6314), .A2(g3934), .ZN(g9634) );
AND2_X4 U_g9635 ( .A1(g6232), .A2(g3937), .ZN(g9635) );
AND4_X4 U_I16735 ( .A1(g5856), .A2(g4338), .A3(g4339), .A4(g5141), .ZN(I16735) );
AND4_X4 U_I16736 ( .A1(g5713), .A2(g5958), .A3(g4735), .A4(g4736), .ZN(I16736) );
AND2_X4 U_g9636 ( .A1(I16735), .A2(I16736), .ZN(g9636) );
AND2_X4 U_g9639 ( .A1(g5438), .A2(g408), .ZN(g9639) );
AND2_X4 U_g9647 ( .A1(g6678), .A2(g3942), .ZN(g9647) );
AND2_X4 U_g9648 ( .A1(g6678), .A2(g3945), .ZN(g9648) );
AND2_X4 U_g9660 ( .A1(g3410), .A2(g3948), .ZN(g9660) );
AND2_X4 U_g9661 ( .A1(g6519), .A2(g3951), .ZN(g9661) );
AND2_X4 U_g9662 ( .A1(g6369), .A2(g3954), .ZN(g9662) );
AND2_X4 U_g9663 ( .A1(g3410), .A2(g3957), .ZN(g9663) );
AND2_X4 U_g9664 ( .A1(g6519), .A2(g3960), .ZN(g9664) );
AND2_X4 U_g9665 ( .A1(g6369), .A2(g3963), .ZN(g9665) );
AND3_X4 U_g9676 ( .A1(g7788), .A2(g6145), .A3(g1224), .ZN(g9676) );
AND2_X4 U_g9722 ( .A1(g3566), .A2(g3966), .ZN(g9722) );
AND2_X4 U_g9723 ( .A1(g6783), .A2(g3969), .ZN(g9723) );
AND2_X4 U_g9724 ( .A1(g6574), .A2(g3972), .ZN(g9724) );
AND2_X4 U_g9725 ( .A1(g6783), .A2(g3975), .ZN(g9725) );
AND2_X4 U_g9726 ( .A1(g6574), .A2(g3978), .ZN(g9726) );
AND2_X4 U_g9745 ( .A1(g3722), .A2(g3981), .ZN(g9745) );
AND2_X4 U_g9746 ( .A1(g7085), .A2(g3984), .ZN(g9746) );
AND2_X4 U_g9747 ( .A1(g6838), .A2(g3987), .ZN(g9747) );
AND2_X4 U_g9748 ( .A1(g6838), .A2(g3990), .ZN(g9748) );
AND2_X4 U_g9759 ( .A1(g3254), .A2(g4000), .ZN(g9759) );
AND2_X4 U_g9760 ( .A1(g6314), .A2(g4003), .ZN(g9760) );
AND2_X4 U_g9761 ( .A1(g6232), .A2(g4006), .ZN(g9761) );
AND2_X4 U_g9762 ( .A1(g3254), .A2(g4009), .ZN(g9762) );
AND2_X4 U_g9763 ( .A1(g6314), .A2(g4012), .ZN(g9763) );
AND2_X4 U_g9764 ( .A1(g6448), .A2(g411), .ZN(g9764) );
AND2_X4 U_g9765 ( .A1(g5438), .A2(g417), .ZN(g9765) );
AND2_X4 U_g9766 ( .A1(g5438), .A2(g4017), .ZN(g9766) );
AND2_X4 U_g9773 ( .A1(g6912), .A2(g4020), .ZN(g9773) );
AND2_X4 U_g9774 ( .A1(g6678), .A2(g4023), .ZN(g9774) );
AND2_X4 U_g9775 ( .A1(g6912), .A2(g4026), .ZN(g9775) );
AND2_X4 U_g9776 ( .A1(g3410), .A2(g4029), .ZN(g9776) );
AND2_X4 U_g9777 ( .A1(g6519), .A2(g4032), .ZN(g9777) );
AND2_X4 U_g9778 ( .A1(g6369), .A2(g4035), .ZN(g9778) );
AND2_X4 U_g9779 ( .A1(g3410), .A2(g4038), .ZN(g9779) );
AND2_X4 U_g9780 ( .A1(g6519), .A2(g4041), .ZN(g9780) );
AND2_X4 U_g9781 ( .A1(g6369), .A2(g4044), .ZN(g9781) );
AND4_X4 U_I16826 ( .A1(g5903), .A2(g4507), .A3(g4508), .A4(g5234), .ZN(I16826) );
AND4_X4 U_I16827 ( .A1(g5771), .A2(g5987), .A3(g4911), .A4(g4912), .ZN(I16827) );
AND2_X4 U_g9782 ( .A1(I16826), .A2(I16827), .ZN(g9782) );
AND2_X4 U_g9785 ( .A1(g5473), .A2(g1095), .ZN(g9785) );
AND2_X4 U_g9793 ( .A1(g6980), .A2(g4049), .ZN(g9793) );
AND2_X4 U_g9794 ( .A1(g6980), .A2(g4052), .ZN(g9794) );
AND2_X4 U_g9806 ( .A1(g3566), .A2(g4055), .ZN(g9806) );
AND2_X4 U_g9807 ( .A1(g6783), .A2(g4058), .ZN(g9807) );
AND2_X4 U_g9808 ( .A1(g6574), .A2(g4061), .ZN(g9808) );
AND2_X4 U_g9809 ( .A1(g3566), .A2(g4064), .ZN(g9809) );
AND2_X4 U_g9810 ( .A1(g6783), .A2(g4067), .ZN(g9810) );
AND2_X4 U_g9811 ( .A1(g6574), .A2(g4070), .ZN(g9811) );
AND3_X4 U_g9822 ( .A1(g7802), .A2(g6166), .A3(g1918), .ZN(g9822) );
AND2_X4 U_g9868 ( .A1(g3722), .A2(g4073), .ZN(g9868) );
AND2_X4 U_g9869 ( .A1(g7085), .A2(g4076), .ZN(g9869) );
AND2_X4 U_g9870 ( .A1(g6838), .A2(g4079), .ZN(g9870) );
AND2_X4 U_g9871 ( .A1(g7085), .A2(g4082), .ZN(g9871) );
AND2_X4 U_g9872 ( .A1(g6838), .A2(g4085), .ZN(g9872) );
AND2_X4 U_g9887 ( .A1(g6232), .A2(g4095), .ZN(g9887) );
AND2_X4 U_g9888 ( .A1(g3254), .A2(g4098), .ZN(g9888) );
AND2_X4 U_g9889 ( .A1(g6314), .A2(g4101), .ZN(g9889) );
AND2_X4 U_g9890 ( .A1(g6232), .A2(g4104), .ZN(g9890) );
AND2_X4 U_g9891 ( .A1(g3254), .A2(g4107), .ZN(g9891) );
AND2_X4 U_g9892 ( .A1(g3306), .A2(g414), .ZN(g9892) );
AND2_X4 U_g9893 ( .A1(g6448), .A2(g420), .ZN(g9893) );
AND2_X4 U_g9894 ( .A1(g6448), .A2(g4112), .ZN(g9894) );
AND2_X4 U_g9901 ( .A1(g3366), .A2(g4115), .ZN(g9901) );
AND2_X4 U_g9902 ( .A1(g6912), .A2(g4118), .ZN(g9902) );
AND2_X4 U_g9903 ( .A1(g6678), .A2(g4121), .ZN(g9903) );
AND2_X4 U_g9904 ( .A1(g3366), .A2(g4124), .ZN(g9904) );
AND2_X4 U_g9905 ( .A1(g3410), .A2(g4127), .ZN(g9905) );
AND2_X4 U_g9906 ( .A1(g6519), .A2(g4130), .ZN(g9906) );
AND2_X4 U_g9907 ( .A1(g6369), .A2(g4133), .ZN(g9907) );
AND2_X4 U_g9908 ( .A1(g3410), .A2(g4136), .ZN(g9908) );
AND2_X4 U_g9909 ( .A1(g6519), .A2(g4139), .ZN(g9909) );
AND2_X4 U_g9910 ( .A1(g6713), .A2(g1098), .ZN(g9910) );
AND2_X4 U_g9911 ( .A1(g5473), .A2(g1104), .ZN(g9911) );
AND2_X4 U_g9912 ( .A1(g5473), .A2(g4144), .ZN(g9912) );
AND2_X4 U_g9919 ( .A1(g7162), .A2(g4147), .ZN(g9919) );
AND2_X4 U_g9920 ( .A1(g6980), .A2(g4150), .ZN(g9920) );
AND2_X4 U_g9921 ( .A1(g7162), .A2(g4153), .ZN(g9921) );
AND2_X4 U_g9922 ( .A1(g3566), .A2(g4156), .ZN(g9922) );
AND2_X4 U_g9923 ( .A1(g6783), .A2(g4159), .ZN(g9923) );
AND2_X4 U_g9924 ( .A1(g6574), .A2(g4162), .ZN(g9924) );
AND2_X4 U_g9925 ( .A1(g3566), .A2(g4165), .ZN(g9925) );
AND2_X4 U_g9926 ( .A1(g6783), .A2(g4168), .ZN(g9926) );
AND2_X4 U_g9927 ( .A1(g6574), .A2(g4171), .ZN(g9927) );
AND4_X4 U_I16930 ( .A1(g5942), .A2(g4683), .A3(g4684), .A4(g5297), .ZN(I16930) );
AND4_X4 U_I16931 ( .A1(g5830), .A2(g6024), .A3(g5070), .A4(g5071), .ZN(I16931) );
AND2_X4 U_g9928 ( .A1(I16930), .A2(I16931), .ZN(g9928) );
AND2_X4 U_g9931 ( .A1(g5512), .A2(g1789), .ZN(g9931) );
AND2_X4 U_g9939 ( .A1(g7230), .A2(g4176), .ZN(g9939) );
AND2_X4 U_g9940 ( .A1(g7230), .A2(g4179), .ZN(g9940) );
AND2_X4 U_g9952 ( .A1(g3722), .A2(g4182), .ZN(g9952) );
AND2_X4 U_g9953 ( .A1(g7085), .A2(g4185), .ZN(g9953) );
AND2_X4 U_g9954 ( .A1(g6838), .A2(g4188), .ZN(g9954) );
AND2_X4 U_g9955 ( .A1(g3722), .A2(g4191), .ZN(g9955) );
AND2_X4 U_g9956 ( .A1(g7085), .A2(g4194), .ZN(g9956) );
AND2_X4 U_g9957 ( .A1(g6838), .A2(g4197), .ZN(g9957) );
AND3_X4 U_g9968 ( .A1(g7815), .A2(g6193), .A3(g2612), .ZN(g9968) );
AND2_X4 U_g10007 ( .A1(g6314), .A2(g4205), .ZN(g10007) );
AND2_X4 U_g10008 ( .A1(g6232), .A2(g4208), .ZN(g10008) );
AND2_X4 U_g10009 ( .A1(g3254), .A2(g4211), .ZN(g10009) );
AND2_X4 U_g10010 ( .A1(g6314), .A2(g4214), .ZN(g10010) );
AND2_X4 U_g10011 ( .A1(g5438), .A2(g4217), .ZN(g10011) );
AND2_X4 U_g10012 ( .A1(g3306), .A2(g423), .ZN(g10012) );
AND2_X4 U_g10013 ( .A1(g3306), .A2(g4221), .ZN(g10013) );
AND2_X4 U_g10014 ( .A1(g5438), .A2(g429), .ZN(g10014) );
AND2_X4 U_g10024 ( .A1(g3398), .A2(g6912), .ZN(g10024) );
AND2_X4 U_g10035 ( .A1(g3366), .A2(g4225), .ZN(g10035) );
AND2_X4 U_g10036 ( .A1(g6912), .A2(g4228), .ZN(g10036) );
AND2_X4 U_g10037 ( .A1(g6678), .A2(g4231), .ZN(g10037) );
AND2_X4 U_g10041 ( .A1(g6369), .A2(g4234), .ZN(g10041) );
AND2_X4 U_g10042 ( .A1(g3410), .A2(g4237), .ZN(g10042) );
AND2_X4 U_g10043 ( .A1(g6519), .A2(g4240), .ZN(g10043) );
AND2_X4 U_g10044 ( .A1(g6369), .A2(g4243), .ZN(g10044) );
AND2_X4 U_g10045 ( .A1(g3410), .A2(g4246), .ZN(g10045) );
AND2_X4 U_g10046 ( .A1(g3462), .A2(g1101), .ZN(g10046) );
AND2_X4 U_g10047 ( .A1(g6713), .A2(g1107), .ZN(g10047) );
AND2_X4 U_g10048 ( .A1(g6713), .A2(g4251), .ZN(g10048) );
AND2_X4 U_g10055 ( .A1(g3522), .A2(g4254), .ZN(g10055) );
AND2_X4 U_g10056 ( .A1(g7162), .A2(g4257), .ZN(g10056) );
AND2_X4 U_g10057 ( .A1(g6980), .A2(g4260), .ZN(g10057) );
AND2_X4 U_g10058 ( .A1(g3522), .A2(g4263), .ZN(g10058) );
AND2_X4 U_g10059 ( .A1(g3566), .A2(g4266), .ZN(g10059) );
AND2_X4 U_g10060 ( .A1(g6783), .A2(g4269), .ZN(g10060) );
AND2_X4 U_g10061 ( .A1(g6574), .A2(g4272), .ZN(g10061) );
AND2_X4 U_g10062 ( .A1(g3566), .A2(g4275), .ZN(g10062) );
AND2_X4 U_g10063 ( .A1(g6783), .A2(g4278), .ZN(g10063) );
AND2_X4 U_g10064 ( .A1(g7015), .A2(g1792), .ZN(g10064) );
AND2_X4 U_g10065 ( .A1(g5512), .A2(g1798), .ZN(g10065) );
AND2_X4 U_g10066 ( .A1(g5512), .A2(g4283), .ZN(g10066) );
AND2_X4 U_g10073 ( .A1(g7358), .A2(g4286), .ZN(g10073) );
AND2_X4 U_g10074 ( .A1(g7230), .A2(g4289), .ZN(g10074) );
AND2_X4 U_g10075 ( .A1(g7358), .A2(g4292), .ZN(g10075) );
AND2_X4 U_g10076 ( .A1(g3722), .A2(g4295), .ZN(g10076) );
AND2_X4 U_g10077 ( .A1(g7085), .A2(g4298), .ZN(g10077) );
AND2_X4 U_g10078 ( .A1(g6838), .A2(g4301), .ZN(g10078) );
AND2_X4 U_g10079 ( .A1(g3722), .A2(g4304), .ZN(g10079) );
AND2_X4 U_g10080 ( .A1(g7085), .A2(g4307), .ZN(g10080) );
AND2_X4 U_g10081 ( .A1(g6838), .A2(g4310), .ZN(g10081) );
AND4_X4 U_I17042 ( .A1(g5976), .A2(g4860), .A3(g4861), .A4(g5334), .ZN(I17042) );
AND4_X4 U_I17043 ( .A1(g5886), .A2(g6040), .A3(g5199), .A4(g5200), .ZN(I17043) );
AND2_X4 U_g10082 ( .A1(I17042), .A2(I17043), .ZN(g10082) );
AND2_X4 U_g10085 ( .A1(g5556), .A2(g2483), .ZN(g10085) );
AND2_X4 U_g10093 ( .A1(g7426), .A2(g4315), .ZN(g10093) );
AND2_X4 U_g10094 ( .A1(g7426), .A2(g4318), .ZN(g10094) );
AND2_X4 U_g10101 ( .A1(g3254), .A2(g4329), .ZN(g10101) );
AND2_X4 U_g10102 ( .A1(g6314), .A2(g4332), .ZN(g10102) );
AND2_X4 U_g10103 ( .A1(g3254), .A2(g4335), .ZN(g10103) );
AND2_X4 U_g10104 ( .A1(g6448), .A2(g4340), .ZN(g10104) );
AND2_X4 U_g10105 ( .A1(g5438), .A2(g4343), .ZN(g10105) );
AND2_X4 U_g10106 ( .A1(g6448), .A2(g432), .ZN(g10106) );
AND2_X4 U_g10107 ( .A1(g5438), .A2(g438), .ZN(g10107) );
AND2_X4 U_g10108 ( .A1(g6486), .A2(g569), .ZN(g10108) );
AND2_X4 U_g10112 ( .A1(g3366), .A2(g4348), .ZN(g10112) );
AND2_X4 U_g10113 ( .A1(g6912), .A2(g4351), .ZN(g10113) );
AND2_X4 U_g10114 ( .A1(g6678), .A2(g4354), .ZN(g10114) );
AND2_X4 U_g10115 ( .A1(g6678), .A2(g4357), .ZN(g10115) );
AND2_X4 U_g10116 ( .A1(g6519), .A2(g4360), .ZN(g10116) );
AND2_X4 U_g10117 ( .A1(g6369), .A2(g4363), .ZN(g10117) );
AND2_X4 U_g10118 ( .A1(g3410), .A2(g4366), .ZN(g10118) );
AND2_X4 U_g10119 ( .A1(g6519), .A2(g4369), .ZN(g10119) );
AND2_X4 U_g10120 ( .A1(g5473), .A2(g4372), .ZN(g10120) );
AND2_X4 U_g10121 ( .A1(g3462), .A2(g1110), .ZN(g10121) );
AND2_X4 U_g10122 ( .A1(g3462), .A2(g4376), .ZN(g10122) );
AND2_X4 U_g10123 ( .A1(g5473), .A2(g1116), .ZN(g10123) );
AND2_X4 U_g10133 ( .A1(g3554), .A2(g7162), .ZN(g10133) );
AND2_X4 U_g10144 ( .A1(g3522), .A2(g4380), .ZN(g10144) );
AND2_X4 U_g10145 ( .A1(g7162), .A2(g4383), .ZN(g10145) );
AND2_X4 U_g10146 ( .A1(g6980), .A2(g4386), .ZN(g10146) );
AND2_X4 U_g10150 ( .A1(g6574), .A2(g4389), .ZN(g10150) );
AND2_X4 U_g10151 ( .A1(g3566), .A2(g4392), .ZN(g10151) );
AND2_X4 U_g10152 ( .A1(g6783), .A2(g4395), .ZN(g10152) );
AND2_X4 U_g10153 ( .A1(g6574), .A2(g4398), .ZN(g10153) );
AND2_X4 U_g10154 ( .A1(g3566), .A2(g4401), .ZN(g10154) );
AND2_X4 U_g10155 ( .A1(g3618), .A2(g1795), .ZN(g10155) );
AND2_X4 U_g10156 ( .A1(g7015), .A2(g1801), .ZN(g10156) );
AND2_X4 U_g10157 ( .A1(g7015), .A2(g4406), .ZN(g10157) );
AND2_X4 U_g10164 ( .A1(g3678), .A2(g4409), .ZN(g10164) );
AND2_X4 U_g10165 ( .A1(g7358), .A2(g4412), .ZN(g10165) );
AND2_X4 U_g10166 ( .A1(g7230), .A2(g4415), .ZN(g10166) );
AND2_X4 U_g10167 ( .A1(g3678), .A2(g4418), .ZN(g10167) );
AND2_X4 U_g10168 ( .A1(g3722), .A2(g4421), .ZN(g10168) );
AND2_X4 U_g10169 ( .A1(g7085), .A2(g4424), .ZN(g10169) );
AND2_X4 U_g10170 ( .A1(g6838), .A2(g4427), .ZN(g10170) );
AND2_X4 U_g10171 ( .A1(g3722), .A2(g4430), .ZN(g10171) );
AND2_X4 U_g10172 ( .A1(g7085), .A2(g4433), .ZN(g10172) );
AND2_X4 U_g10173 ( .A1(g7265), .A2(g2486), .ZN(g10173) );
AND2_X4 U_g10174 ( .A1(g5556), .A2(g2492), .ZN(g10174) );
AND2_X4 U_g10175 ( .A1(g5556), .A2(g4438), .ZN(g10175) );
AND2_X4 U_g10182 ( .A1(g7488), .A2(g4441), .ZN(g10182) );
AND2_X4 U_g10183 ( .A1(g7426), .A2(g4444), .ZN(g10183) );
AND2_X4 U_g10184 ( .A1(g7488), .A2(g4447), .ZN(g10184) );
AND4_X4 U_I17156 ( .A1(g6898), .A2(g2998), .A3(g6901), .A4(g3002), .ZN(I17156) );
AND4_X4 U_g10186 ( .A1(g3013), .A2(g7466), .A3(g3024), .A4(I17156), .ZN(g10186) );
AND2_X4 U_g10192 ( .A1(g3254), .A2(g4453), .ZN(g10192) );
AND2_X4 U_g10193 ( .A1(g3306), .A2(g4465), .ZN(g10193) );
AND2_X4 U_g10194 ( .A1(g6448), .A2(g4468), .ZN(g10194) );
AND2_X4 U_g10195 ( .A1(g5438), .A2(g4471), .ZN(g10195) );
AND2_X4 U_g10196 ( .A1(g3306), .A2(g435), .ZN(g10196) );
AND2_X4 U_g10197 ( .A1(g6448), .A2(g441), .ZN(g10197) );
AND2_X4 U_g10198 ( .A1(g6643), .A2(g571), .ZN(g10198) );
AND2_X4 U_g10199 ( .A1(g6486), .A2(g4476), .ZN(g10199) );
AND2_X4 U_g10200 ( .A1(g6486), .A2(g587), .ZN(g10200) );
AND2_X4 U_g10201 ( .A1(g3366), .A2(g4480), .ZN(g10201) );
AND2_X4 U_g10202 ( .A1(g6912), .A2(g4483), .ZN(g10202) );
AND2_X4 U_g10203 ( .A1(g6678), .A2(g4486), .ZN(g10203) );
AND2_X4 U_g10204 ( .A1(g6912), .A2(g4489), .ZN(g10204) );
AND2_X4 U_g10205 ( .A1(g6678), .A2(g4492), .ZN(g10205) );
AND2_X4 U_g10206 ( .A1(g3410), .A2(g4498), .ZN(g10206) );
AND2_X4 U_g10207 ( .A1(g6519), .A2(g4501), .ZN(g10207) );
AND2_X4 U_g10208 ( .A1(g3410), .A2(g4504), .ZN(g10208) );
AND2_X4 U_g10209 ( .A1(g6713), .A2(g4509), .ZN(g10209) );
AND2_X4 U_g10210 ( .A1(g5473), .A2(g4512), .ZN(g10210) );
AND2_X4 U_g10211 ( .A1(g6713), .A2(g1119), .ZN(g10211) );
AND2_X4 U_g10212 ( .A1(g5473), .A2(g1125), .ZN(g10212) );
AND2_X4 U_g10213 ( .A1(g6751), .A2(g1255), .ZN(g10213) );
AND2_X4 U_g10217 ( .A1(g3522), .A2(g4517), .ZN(g10217) );
AND2_X4 U_g10218 ( .A1(g7162), .A2(g4520), .ZN(g10218) );
AND2_X4 U_g10219 ( .A1(g6980), .A2(g4523), .ZN(g10219) );
AND2_X4 U_g10220 ( .A1(g6980), .A2(g4526), .ZN(g10220) );
AND2_X4 U_g10221 ( .A1(g6783), .A2(g4529), .ZN(g10221) );
AND2_X4 U_g10222 ( .A1(g6574), .A2(g4532), .ZN(g10222) );
AND2_X4 U_g10223 ( .A1(g3566), .A2(g4535), .ZN(g10223) );
AND2_X4 U_g10224 ( .A1(g6783), .A2(g4538), .ZN(g10224) );
AND2_X4 U_g10225 ( .A1(g5512), .A2(g4541), .ZN(g10225) );
AND2_X4 U_g10226 ( .A1(g3618), .A2(g1804), .ZN(g10226) );
AND2_X4 U_g10227 ( .A1(g3618), .A2(g4545), .ZN(g10227) );
AND2_X4 U_g10228 ( .A1(g5512), .A2(g1810), .ZN(g10228) );
AND2_X4 U_g10238 ( .A1(g3710), .A2(g7358), .ZN(g10238) );
AND2_X4 U_g10249 ( .A1(g3678), .A2(g4549), .ZN(g10249) );
AND2_X4 U_g10250 ( .A1(g7358), .A2(g4552), .ZN(g10250) );
AND2_X4 U_g10251 ( .A1(g7230), .A2(g4555), .ZN(g10251) );
AND2_X4 U_g10255 ( .A1(g6838), .A2(g4558), .ZN(g10255) );
AND2_X4 U_g10256 ( .A1(g3722), .A2(g4561), .ZN(g10256) );
AND2_X4 U_g10257 ( .A1(g7085), .A2(g4564), .ZN(g10257) );
AND2_X4 U_g10258 ( .A1(g6838), .A2(g4567), .ZN(g10258) );
AND2_X4 U_g10259 ( .A1(g3722), .A2(g4570), .ZN(g10259) );
AND2_X4 U_g10260 ( .A1(g3774), .A2(g2489), .ZN(g10260) );
AND2_X4 U_g10261 ( .A1(g7265), .A2(g2495), .ZN(g10261) );
AND2_X4 U_g10262 ( .A1(g7265), .A2(g4575), .ZN(g10262) );
AND2_X4 U_g10269 ( .A1(g3834), .A2(g4578), .ZN(g10269) );
AND2_X4 U_g10270 ( .A1(g7488), .A2(g4581), .ZN(g10270) );
AND2_X4 U_g10271 ( .A1(g7426), .A2(g4584), .ZN(g10271) );
AND2_X4 U_g10272 ( .A1(g3834), .A2(g4587), .ZN(g10272) );
AND2_X4 U_g10279 ( .A1(g3306), .A2(g4592), .ZN(g10279) );
AND2_X4 U_g10280 ( .A1(g6448), .A2(g4595), .ZN(g10280) );
AND2_X4 U_g10281 ( .A1(g5438), .A2(g4598), .ZN(g10281) );
AND2_X4 U_g10282 ( .A1(g3306), .A2(g444), .ZN(g10282) );
AND2_X4 U_g10283 ( .A1(g3338), .A2(g573), .ZN(g10283) );
AND2_X4 U_g10284 ( .A1(g6643), .A2(g4603), .ZN(g10284) );
AND2_X4 U_g10285 ( .A1(g6486), .A2(g4606), .ZN(g10285) );
AND2_X4 U_g10286 ( .A1(g6643), .A2(g590), .ZN(g10286) );
AND2_X4 U_g10287 ( .A1(g6486), .A2(g596), .ZN(g10287) );
AND2_X4 U_g10288 ( .A1(g3366), .A2(g4611), .ZN(g10288) );
AND2_X4 U_g10289 ( .A1(g6912), .A2(g4614), .ZN(g10289) );
AND2_X4 U_g10290 ( .A1(g6678), .A2(g4617), .ZN(g10290) );
AND2_X4 U_g10291 ( .A1(g3366), .A2(g4620), .ZN(g10291) );
AND2_X4 U_g10292 ( .A1(g6912), .A2(g4623), .ZN(g10292) );
AND2_X4 U_g10293 ( .A1(g6678), .A2(g4626), .ZN(g10293) );
AND2_X4 U_g10294 ( .A1(g3410), .A2(g4629), .ZN(g10294) );
AND2_X4 U_g10295 ( .A1(g3462), .A2(g4641), .ZN(g10295) );
AND2_X4 U_g10296 ( .A1(g6713), .A2(g4644), .ZN(g10296) );
AND2_X4 U_g10297 ( .A1(g5473), .A2(g4647), .ZN(g10297) );
AND2_X4 U_g10298 ( .A1(g3462), .A2(g1122), .ZN(g10298) );
AND2_X4 U_g10299 ( .A1(g6713), .A2(g1128), .ZN(g10299) );
AND2_X4 U_g10300 ( .A1(g6945), .A2(g1257), .ZN(g10300) );
AND2_X4 U_g10301 ( .A1(g6751), .A2(g4652), .ZN(g10301) );
AND2_X4 U_g10302 ( .A1(g6751), .A2(g1273), .ZN(g10302) );
AND2_X4 U_g10303 ( .A1(g3522), .A2(g4656), .ZN(g10303) );
AND2_X4 U_g10304 ( .A1(g7162), .A2(g4659), .ZN(g10304) );
AND2_X4 U_g10305 ( .A1(g6980), .A2(g4662), .ZN(g10305) );
AND2_X4 U_g10306 ( .A1(g7162), .A2(g4665), .ZN(g10306) );
AND2_X4 U_g10307 ( .A1(g6980), .A2(g4668), .ZN(g10307) );
AND2_X4 U_g10308 ( .A1(g3566), .A2(g4674), .ZN(g10308) );
AND2_X4 U_g10309 ( .A1(g6783), .A2(g4677), .ZN(g10309) );
AND2_X4 U_g10310 ( .A1(g3566), .A2(g4680), .ZN(g10310) );
AND2_X4 U_g10311 ( .A1(g7015), .A2(g4685), .ZN(g10311) );
AND2_X4 U_g10312 ( .A1(g5512), .A2(g4688), .ZN(g10312) );
AND2_X4 U_g10313 ( .A1(g7015), .A2(g1813), .ZN(g10313) );
AND2_X4 U_g10314 ( .A1(g5512), .A2(g1819), .ZN(g10314) );
AND2_X4 U_g10315 ( .A1(g7053), .A2(g1949), .ZN(g10315) );
AND2_X4 U_g10319 ( .A1(g3678), .A2(g4693), .ZN(g10319) );
AND2_X4 U_g10320 ( .A1(g7358), .A2(g4696), .ZN(g10320) );
AND2_X4 U_g10321 ( .A1(g7230), .A2(g4699), .ZN(g10321) );
AND2_X4 U_g10322 ( .A1(g7230), .A2(g4702), .ZN(g10322) );
AND2_X4 U_g10323 ( .A1(g7085), .A2(g4705), .ZN(g10323) );
AND2_X4 U_g10324 ( .A1(g6838), .A2(g4708), .ZN(g10324) );
AND2_X4 U_g10325 ( .A1(g3722), .A2(g4711), .ZN(g10325) );
AND2_X4 U_g10326 ( .A1(g7085), .A2(g4714), .ZN(g10326) );
AND2_X4 U_g10327 ( .A1(g5556), .A2(g4717), .ZN(g10327) );
AND2_X4 U_g10328 ( .A1(g3774), .A2(g2498), .ZN(g10328) );
AND2_X4 U_g10329 ( .A1(g3774), .A2(g4721), .ZN(g10329) );
AND2_X4 U_g10330 ( .A1(g5556), .A2(g2504), .ZN(g10330) );
AND2_X4 U_g10340 ( .A1(g3866), .A2(g7488), .ZN(g10340) );
AND2_X4 U_g10351 ( .A1(g3834), .A2(g4725), .ZN(g10351) );
AND2_X4 U_g10352 ( .A1(g7488), .A2(g4728), .ZN(g10352) );
AND2_X4 U_g10353 ( .A1(g7426), .A2(g4731), .ZN(g10353) );
AND2_X4 U_g10360 ( .A1(g3306), .A2(g4737), .ZN(g10360) );
AND2_X4 U_g10361 ( .A1(g6448), .A2(g4740), .ZN(g10361) );
AND2_X4 U_g10362 ( .A1(g3338), .A2(g4743), .ZN(g10362) );
AND2_X4 U_g10363 ( .A1(g6643), .A2(g4746), .ZN(g10363) );
AND2_X4 U_g10364 ( .A1(g6486), .A2(g4749), .ZN(g10364) );
AND2_X4 U_g10365 ( .A1(g3338), .A2(g593), .ZN(g10365) );
AND2_X4 U_g10366 ( .A1(g6643), .A2(g599), .ZN(g10366) );
AND2_X4 U_g10367 ( .A1(g3366), .A2(g4754), .ZN(g10367) );
AND2_X4 U_g10368 ( .A1(g6912), .A2(g4757), .ZN(g10368) );
AND2_X4 U_g10369 ( .A1(g6678), .A2(g4760), .ZN(g10369) );
AND2_X4 U_g10370 ( .A1(g3366), .A2(g4763), .ZN(g10370) );
AND2_X4 U_g10371 ( .A1(g6912), .A2(g4766), .ZN(g10371) );
AND2_X4 U_g10372 ( .A1(g3462), .A2(g4769), .ZN(g10372) );
AND2_X4 U_g10373 ( .A1(g6713), .A2(g4772), .ZN(g10373) );
AND2_X4 U_g10374 ( .A1(g5473), .A2(g4775), .ZN(g10374) );
AND2_X4 U_g10375 ( .A1(g3462), .A2(g1131), .ZN(g10375) );
AND2_X4 U_g10376 ( .A1(g3494), .A2(g1259), .ZN(g10376) );
AND2_X4 U_g10377 ( .A1(g6945), .A2(g4780), .ZN(g10377) );
AND2_X4 U_g10378 ( .A1(g6751), .A2(g4783), .ZN(g10378) );
AND2_X4 U_g10379 ( .A1(g6945), .A2(g1276), .ZN(g10379) );
AND2_X4 U_g10380 ( .A1(g6751), .A2(g1282), .ZN(g10380) );
AND2_X4 U_g10381 ( .A1(g3522), .A2(g4788), .ZN(g10381) );
AND2_X4 U_g10382 ( .A1(g7162), .A2(g4791), .ZN(g10382) );
AND2_X4 U_g10383 ( .A1(g6980), .A2(g4794), .ZN(g10383) );
AND2_X4 U_g10384 ( .A1(g3522), .A2(g4797), .ZN(g10384) );
AND2_X4 U_g10385 ( .A1(g7162), .A2(g4800), .ZN(g10385) );
AND2_X4 U_g10386 ( .A1(g6980), .A2(g4803), .ZN(g10386) );
AND2_X4 U_g10387 ( .A1(g3566), .A2(g4806), .ZN(g10387) );
AND2_X4 U_g10388 ( .A1(g3618), .A2(g4818), .ZN(g10388) );
AND2_X4 U_g10389 ( .A1(g7015), .A2(g4821), .ZN(g10389) );
AND2_X4 U_g10390 ( .A1(g5512), .A2(g4824), .ZN(g10390) );
AND2_X4 U_g10391 ( .A1(g3618), .A2(g1816), .ZN(g10391) );
AND2_X4 U_g10392 ( .A1(g7015), .A2(g1822), .ZN(g10392) );
AND2_X4 U_g10393 ( .A1(g7195), .A2(g1951), .ZN(g10393) );
AND2_X4 U_g10394 ( .A1(g7053), .A2(g4829), .ZN(g10394) );
AND2_X4 U_g10395 ( .A1(g7053), .A2(g1967), .ZN(g10395) );
AND2_X4 U_g10396 ( .A1(g3678), .A2(g4833), .ZN(g10396) );
AND2_X4 U_g10397 ( .A1(g7358), .A2(g4836), .ZN(g10397) );
AND2_X4 U_g10398 ( .A1(g7230), .A2(g4839), .ZN(g10398) );
AND2_X4 U_g10399 ( .A1(g7358), .A2(g4842), .ZN(g10399) );
AND2_X4 U_g10400 ( .A1(g7230), .A2(g4845), .ZN(g10400) );
AND2_X4 U_g10401 ( .A1(g3722), .A2(g4851), .ZN(g10401) );
AND2_X4 U_g10402 ( .A1(g7085), .A2(g4854), .ZN(g10402) );
AND2_X4 U_g10403 ( .A1(g3722), .A2(g4857), .ZN(g10403) );
AND2_X4 U_g10404 ( .A1(g7265), .A2(g4862), .ZN(g10404) );
AND2_X4 U_g10405 ( .A1(g5556), .A2(g4865), .ZN(g10405) );
AND2_X4 U_g10406 ( .A1(g7265), .A2(g2507), .ZN(g10406) );
AND2_X4 U_g10407 ( .A1(g5556), .A2(g2513), .ZN(g10407) );
AND2_X4 U_g10408 ( .A1(g7303), .A2(g2643), .ZN(g10408) );
AND2_X4 U_g10412 ( .A1(g3834), .A2(g4870), .ZN(g10412) );
AND2_X4 U_g10413 ( .A1(g7488), .A2(g4873), .ZN(g10413) );
AND2_X4 U_g10414 ( .A1(g7426), .A2(g4876), .ZN(g10414) );
AND2_X4 U_g10415 ( .A1(g7426), .A2(g4879), .ZN(g10415) );
AND2_X4 U_g10422 ( .A1(g3306), .A2(g4882), .ZN(g10422) );
AND2_X4 U_g10423 ( .A1(g5438), .A2(g4885), .ZN(g10423) );
AND2_X4 U_g10430 ( .A1(g3338), .A2(g4888), .ZN(g10430) );
AND2_X4 U_g10431 ( .A1(g6643), .A2(g4891), .ZN(g10431) );
AND2_X4 U_g10432 ( .A1(g6486), .A2(g4894), .ZN(g10432) );
AND2_X4 U_g10433 ( .A1(g3338), .A2(g602), .ZN(g10433) );
AND2_X4 U_g10434 ( .A1(g6486), .A2(g605), .ZN(g10434) );
AND2_X4 U_g10435 ( .A1(g3366), .A2(g4899), .ZN(g10435) );
AND2_X4 U_g10436 ( .A1(g6912), .A2(g4902), .ZN(g10436) );
AND2_X4 U_g10437 ( .A1(g6678), .A2(g4905), .ZN(g10437) );
AND2_X4 U_g10438 ( .A1(g3366), .A2(g4908), .ZN(g10438) );
AND2_X4 U_g10439 ( .A1(g3462), .A2(g4913), .ZN(g10439) );
AND2_X4 U_g10440 ( .A1(g6713), .A2(g4916), .ZN(g10440) );
AND2_X4 U_g10441 ( .A1(g3494), .A2(g4919), .ZN(g10441) );
AND2_X4 U_g10442 ( .A1(g6945), .A2(g4922), .ZN(g10442) );
AND2_X4 U_g10443 ( .A1(g6751), .A2(g4925), .ZN(g10443) );
AND2_X4 U_g10444 ( .A1(g3494), .A2(g1279), .ZN(g10444) );
AND2_X4 U_g10445 ( .A1(g6945), .A2(g1285), .ZN(g10445) );
AND2_X4 U_g10446 ( .A1(g3522), .A2(g4930), .ZN(g10446) );
AND2_X4 U_g10447 ( .A1(g7162), .A2(g4933), .ZN(g10447) );
AND2_X4 U_g10448 ( .A1(g6980), .A2(g4936), .ZN(g10448) );
AND2_X4 U_g10449 ( .A1(g3522), .A2(g4939), .ZN(g10449) );
AND2_X4 U_g10450 ( .A1(g7162), .A2(g4942), .ZN(g10450) );
AND2_X4 U_g10451 ( .A1(g3618), .A2(g4945), .ZN(g10451) );
AND2_X4 U_g10452 ( .A1(g7015), .A2(g4948), .ZN(g10452) );
AND2_X4 U_g10453 ( .A1(g5512), .A2(g4951), .ZN(g10453) );
AND2_X4 U_g10454 ( .A1(g3618), .A2(g1825), .ZN(g10454) );
AND2_X4 U_g10455 ( .A1(g3650), .A2(g1953), .ZN(g10455) );
AND2_X4 U_g10456 ( .A1(g7195), .A2(g4956), .ZN(g10456) );
AND2_X4 U_g10457 ( .A1(g7053), .A2(g4959), .ZN(g10457) );
AND2_X4 U_g10458 ( .A1(g7195), .A2(g1970), .ZN(g10458) );
AND2_X4 U_g10459 ( .A1(g7053), .A2(g1976), .ZN(g10459) );
AND2_X4 U_g10460 ( .A1(g3678), .A2(g4964), .ZN(g10460) );
AND2_X4 U_g10461 ( .A1(g7358), .A2(g4967), .ZN(g10461) );
AND2_X4 U_g10462 ( .A1(g7230), .A2(g4970), .ZN(g10462) );
AND2_X4 U_g10463 ( .A1(g3678), .A2(g4973), .ZN(g10463) );
AND2_X4 U_g10464 ( .A1(g7358), .A2(g4976), .ZN(g10464) );
AND2_X4 U_g10465 ( .A1(g7230), .A2(g4979), .ZN(g10465) );
AND2_X4 U_g10466 ( .A1(g3722), .A2(g4982), .ZN(g10466) );
AND2_X4 U_g10467 ( .A1(g3774), .A2(g4994), .ZN(g10467) );
AND2_X4 U_g10468 ( .A1(g7265), .A2(g4997), .ZN(g10468) );
AND2_X4 U_g10469 ( .A1(g5556), .A2(g5000), .ZN(g10469) );
AND2_X4 U_g10470 ( .A1(g3774), .A2(g2510), .ZN(g10470) );
AND2_X4 U_g10471 ( .A1(g7265), .A2(g2516), .ZN(g10471) );
AND2_X4 U_g10472 ( .A1(g7391), .A2(g2645), .ZN(g10472) );
AND2_X4 U_g10473 ( .A1(g7303), .A2(g5005), .ZN(g10473) );
AND2_X4 U_g10474 ( .A1(g7303), .A2(g2661), .ZN(g10474) );
AND2_X4 U_g10475 ( .A1(g3834), .A2(g5009), .ZN(g10475) );
AND2_X4 U_g10476 ( .A1(g7488), .A2(g5012), .ZN(g10476) );
AND2_X4 U_g10477 ( .A1(g7426), .A2(g5015), .ZN(g10477) );
AND2_X4 U_g10478 ( .A1(g7488), .A2(g5018), .ZN(g10478) );
AND2_X4 U_g10479 ( .A1(g7426), .A2(g5021), .ZN(g10479) );
AND3_X4 U_I17429 ( .A1(g6901), .A2(g7338), .A3(g7146), .ZN(I17429) );
AND3_X4 U_g10480 ( .A1(g7466), .A2(g7342), .A3(I17429), .ZN(g10480) );
AND2_X4 U_g10485 ( .A1(g6448), .A2(g5024), .ZN(g10485) );
AND2_X4 U_g10492 ( .A1(g3338), .A2(g5027), .ZN(g10492) );
AND2_X4 U_g10493 ( .A1(g6643), .A2(g5030), .ZN(g10493) );
AND2_X4 U_g10494 ( .A1(g6643), .A2(g608), .ZN(g10494) );
AND2_X4 U_g10495 ( .A1(g6486), .A2(g614), .ZN(g10495) );
AND2_X4 U_g10496 ( .A1(g3366), .A2(g5035), .ZN(g10496) );
AND2_X4 U_g10497 ( .A1(g6912), .A2(g5038), .ZN(g10497) );
AND2_X4 U_g10498 ( .A1(g3462), .A2(g5041), .ZN(g10498) );
AND2_X4 U_g10499 ( .A1(g5473), .A2(g5044), .ZN(g10499) );
AND2_X4 U_g10506 ( .A1(g3494), .A2(g5047), .ZN(g10506) );
AND2_X4 U_g10507 ( .A1(g6945), .A2(g5050), .ZN(g10507) );
AND2_X4 U_g10508 ( .A1(g6751), .A2(g5053), .ZN(g10508) );
AND2_X4 U_g10509 ( .A1(g3494), .A2(g1288), .ZN(g10509) );
AND2_X4 U_g10510 ( .A1(g6751), .A2(g1291), .ZN(g10510) );
AND2_X4 U_g10511 ( .A1(g3522), .A2(g5058), .ZN(g10511) );
AND2_X4 U_g10512 ( .A1(g7162), .A2(g5061), .ZN(g10512) );
AND2_X4 U_g10513 ( .A1(g6980), .A2(g5064), .ZN(g10513) );
AND2_X4 U_g10514 ( .A1(g3522), .A2(g5067), .ZN(g10514) );
AND2_X4 U_g10515 ( .A1(g3618), .A2(g5072), .ZN(g10515) );
AND2_X4 U_g10516 ( .A1(g7015), .A2(g5075), .ZN(g10516) );
AND2_X4 U_g10517 ( .A1(g3650), .A2(g5078), .ZN(g10517) );
AND2_X4 U_g10518 ( .A1(g7195), .A2(g5081), .ZN(g10518) );
AND2_X4 U_g10519 ( .A1(g7053), .A2(g5084), .ZN(g10519) );
AND2_X4 U_g10520 ( .A1(g3650), .A2(g1973), .ZN(g10520) );
AND2_X4 U_g10521 ( .A1(g7195), .A2(g1979), .ZN(g10521) );
AND2_X4 U_g10522 ( .A1(g3678), .A2(g5089), .ZN(g10522) );
AND2_X4 U_g10523 ( .A1(g7358), .A2(g5092), .ZN(g10523) );
AND2_X4 U_g10524 ( .A1(g7230), .A2(g5095), .ZN(g10524) );
AND2_X4 U_g10525 ( .A1(g3678), .A2(g5098), .ZN(g10525) );
AND2_X4 U_g10526 ( .A1(g7358), .A2(g5101), .ZN(g10526) );
AND2_X4 U_g10527 ( .A1(g3774), .A2(g5104), .ZN(g10527) );
AND2_X4 U_g10528 ( .A1(g7265), .A2(g5107), .ZN(g10528) );
AND2_X4 U_g10529 ( .A1(g5556), .A2(g5110), .ZN(g10529) );
AND2_X4 U_g10530 ( .A1(g3774), .A2(g2519), .ZN(g10530) );
AND2_X4 U_g10531 ( .A1(g3806), .A2(g2647), .ZN(g10531) );
AND2_X4 U_g10532 ( .A1(g7391), .A2(g5115), .ZN(g10532) );
AND2_X4 U_g10533 ( .A1(g7303), .A2(g5118), .ZN(g10533) );
AND2_X4 U_g10534 ( .A1(g7391), .A2(g2664), .ZN(g10534) );
AND2_X4 U_g10535 ( .A1(g7303), .A2(g2670), .ZN(g10535) );
AND2_X4 U_g10536 ( .A1(g3834), .A2(g5123), .ZN(g10536) );
AND2_X4 U_g10537 ( .A1(g7488), .A2(g5126), .ZN(g10537) );
AND2_X4 U_g10538 ( .A1(g7426), .A2(g5129), .ZN(g10538) );
AND2_X4 U_g10539 ( .A1(g3834), .A2(g5132), .ZN(g10539) );
AND2_X4 U_g10540 ( .A1(g7488), .A2(g5135), .ZN(g10540) );
AND2_X4 U_g10541 ( .A1(g7426), .A2(g5138), .ZN(g10541) );
AND2_X4 U_g10548 ( .A1(g3306), .A2(g5142), .ZN(g10548) );
AND2_X4 U_g10555 ( .A1(g3338), .A2(g5145), .ZN(g10555) );
AND2_X4 U_g10556 ( .A1(g3338), .A2(g611), .ZN(g10556) );
AND2_X4 U_g10557 ( .A1(g6643), .A2(g617), .ZN(g10557) );
AND2_X4 U_g10558 ( .A1(g3366), .A2(g5150), .ZN(g10558) );
AND2_X4 U_g10559 ( .A1(g6713), .A2(g5153), .ZN(g10559) );
AND2_X4 U_g10566 ( .A1(g3494), .A2(g5156), .ZN(g10566) );
AND2_X4 U_g10567 ( .A1(g6945), .A2(g5159), .ZN(g10567) );
AND2_X4 U_g10568 ( .A1(g6945), .A2(g1294), .ZN(g10568) );
AND2_X4 U_g10569 ( .A1(g6751), .A2(g1300), .ZN(g10569) );
AND2_X4 U_g10570 ( .A1(g3522), .A2(g5164), .ZN(g10570) );
AND2_X4 U_g10571 ( .A1(g7162), .A2(g5167), .ZN(g10571) );
AND2_X4 U_g10572 ( .A1(g3618), .A2(g5170), .ZN(g10572) );
AND2_X4 U_g10573 ( .A1(g5512), .A2(g5173), .ZN(g10573) );
AND2_X4 U_g10580 ( .A1(g3650), .A2(g5176), .ZN(g10580) );
AND2_X4 U_g10581 ( .A1(g7195), .A2(g5179), .ZN(g10581) );
AND2_X4 U_g10582 ( .A1(g7053), .A2(g5182), .ZN(g10582) );
AND2_X4 U_g10583 ( .A1(g3650), .A2(g1982), .ZN(g10583) );
AND2_X4 U_g10584 ( .A1(g7053), .A2(g1985), .ZN(g10584) );
AND2_X4 U_g10585 ( .A1(g3678), .A2(g5187), .ZN(g10585) );
AND2_X4 U_g10586 ( .A1(g7358), .A2(g5190), .ZN(g10586) );
AND2_X4 U_g10587 ( .A1(g7230), .A2(g5193), .ZN(g10587) );
AND2_X4 U_g10588 ( .A1(g3678), .A2(g5196), .ZN(g10588) );
AND2_X4 U_g10589 ( .A1(g3774), .A2(g5201), .ZN(g10589) );
AND2_X4 U_g10590 ( .A1(g7265), .A2(g5204), .ZN(g10590) );
AND2_X4 U_g10591 ( .A1(g3806), .A2(g5207), .ZN(g10591) );
AND2_X4 U_g10592 ( .A1(g7391), .A2(g5210), .ZN(g10592) );
AND2_X4 U_g10593 ( .A1(g7303), .A2(g5213), .ZN(g10593) );
AND2_X4 U_g10594 ( .A1(g3806), .A2(g2667), .ZN(g10594) );
AND2_X4 U_g10595 ( .A1(g7391), .A2(g2673), .ZN(g10595) );
AND2_X4 U_g10596 ( .A1(g3834), .A2(g5218), .ZN(g10596) );
AND2_X4 U_g10597 ( .A1(g7488), .A2(g5221), .ZN(g10597) );
AND2_X4 U_g10598 ( .A1(g7426), .A2(g5224), .ZN(g10598) );
AND2_X4 U_g10599 ( .A1(g3834), .A2(g5227), .ZN(g10599) );
AND2_X4 U_g10600 ( .A1(g7488), .A2(g5230), .ZN(g10600) );
AND2_X4 U_g10604 ( .A1(g3338), .A2(g620), .ZN(g10604) );
AND2_X4 U_g10605 ( .A1(g3462), .A2(g5235), .ZN(g10605) );
AND2_X4 U_g10612 ( .A1(g3494), .A2(g5238), .ZN(g10612) );
AND2_X4 U_g10613 ( .A1(g3494), .A2(g1297), .ZN(g10613) );
AND2_X4 U_g10614 ( .A1(g6945), .A2(g1303), .ZN(g10614) );
AND2_X4 U_g10615 ( .A1(g3522), .A2(g5243), .ZN(g10615) );
AND2_X4 U_g10616 ( .A1(g7015), .A2(g5246), .ZN(g10616) );
AND2_X4 U_g10623 ( .A1(g3650), .A2(g5249), .ZN(g10623) );
AND2_X4 U_g10624 ( .A1(g7195), .A2(g5252), .ZN(g10624) );
AND2_X4 U_g10625 ( .A1(g7195), .A2(g1988), .ZN(g10625) );
AND2_X4 U_g10626 ( .A1(g7053), .A2(g1994), .ZN(g10626) );
AND2_X4 U_g10627 ( .A1(g3678), .A2(g5257), .ZN(g10627) );
AND2_X4 U_g10628 ( .A1(g7358), .A2(g5260), .ZN(g10628) );
AND2_X4 U_g10629 ( .A1(g3774), .A2(g5263), .ZN(g10629) );
AND2_X4 U_g10630 ( .A1(g5556), .A2(g5266), .ZN(g10630) );
AND2_X4 U_g10637 ( .A1(g3806), .A2(g5269), .ZN(g10637) );
AND2_X4 U_g10638 ( .A1(g7391), .A2(g5272), .ZN(g10638) );
AND2_X4 U_g10639 ( .A1(g7303), .A2(g5275), .ZN(g10639) );
AND2_X4 U_g10640 ( .A1(g3806), .A2(g2676), .ZN(g10640) );
AND2_X4 U_g10641 ( .A1(g7303), .A2(g2679), .ZN(g10641) );
AND2_X4 U_g10642 ( .A1(g3834), .A2(g5280), .ZN(g10642) );
AND2_X4 U_g10643 ( .A1(g7488), .A2(g5283), .ZN(g10643) );
AND2_X4 U_g10644 ( .A1(g7426), .A2(g5286), .ZN(g10644) );
AND2_X4 U_g10645 ( .A1(g3834), .A2(g5289), .ZN(g10645) );
AND2_X4 U_g10650 ( .A1(g6678), .A2(g5293), .ZN(g10650) );
AND2_X4 U_g10651 ( .A1(g3494), .A2(g1306), .ZN(g10651) );
AND2_X4 U_g10652 ( .A1(g3618), .A2(g5298), .ZN(g10652) );
AND2_X4 U_g10659 ( .A1(g3650), .A2(g5301), .ZN(g10659) );
AND2_X4 U_g10660 ( .A1(g3650), .A2(g1991), .ZN(g10660) );
AND2_X4 U_g10661 ( .A1(g7195), .A2(g1997), .ZN(g10661) );
AND2_X4 U_g10662 ( .A1(g3678), .A2(g5306), .ZN(g10662) );
AND2_X4 U_g10663 ( .A1(g7265), .A2(g5309), .ZN(g10663) );
AND2_X4 U_g10670 ( .A1(g3806), .A2(g5312), .ZN(g10670) );
AND2_X4 U_g10671 ( .A1(g7391), .A2(g5315), .ZN(g10671) );
AND2_X4 U_g10672 ( .A1(g7391), .A2(g2682), .ZN(g10672) );
AND2_X4 U_g10673 ( .A1(g7303), .A2(g2688), .ZN(g10673) );
AND2_X4 U_g10674 ( .A1(g3834), .A2(g5320), .ZN(g10674) );
AND2_X4 U_g10675 ( .A1(g7488), .A2(g5323), .ZN(g10675) );
AND2_X4 U_g10678 ( .A1(g6912), .A2(g5327), .ZN(g10678) );
AND2_X4 U_g10680 ( .A1(g6980), .A2(g5330), .ZN(g10680) );
AND2_X4 U_g10681 ( .A1(g3650), .A2(g2000), .ZN(g10681) );
AND2_X4 U_g10682 ( .A1(g3774), .A2(g5335), .ZN(g10682) );
AND2_X4 U_g10689 ( .A1(g3806), .A2(g5338), .ZN(g10689) );
AND2_X4 U_g10690 ( .A1(g3806), .A2(g2685), .ZN(g10690) );
AND2_X4 U_g10691 ( .A1(g7391), .A2(g2691), .ZN(g10691) );
AND2_X4 U_g10692 ( .A1(g3834), .A2(g5343), .ZN(g10692) );
AND4_X4 U_g10693 ( .A1(g7462), .A2(g7522), .A3(g2924), .A4(g7545), .ZN(g10693) );
AND2_X4 U_g10704 ( .A1(g3366), .A2(g5352), .ZN(g10704) );
AND2_X4 U_g10707 ( .A1(g7162), .A2(g5355), .ZN(g10707) );
AND2_X4 U_g10709 ( .A1(g7230), .A2(g5358), .ZN(g10709) );
AND2_X4 U_g10710 ( .A1(g3806), .A2(g2694), .ZN(g10710) );
AND3_X4 U_I17599 ( .A1(g7566), .A2(g7583), .A3(g7587), .ZN(I17599) );
AND3_X4 U_g10711 ( .A1(g7595), .A2(g7600), .A3(I17599), .ZN(g10711) );
AND2_X4 U_g10724 ( .A1(g3522), .A2(g5369), .ZN(g10724) );
AND2_X4 U_g10727 ( .A1(g7358), .A2(g5372), .ZN(g10727) );
AND2_X4 U_g10729 ( .A1(g7426), .A2(g5375), .ZN(g10729) );
AND2_X4 U_g10745 ( .A1(g3678), .A2(g5382), .ZN(g10745) );
AND2_X4 U_g10748 ( .A1(g7488), .A2(g5385), .ZN(g10748) );
AND2_X4 U_g10764 ( .A1(g3834), .A2(g5391), .ZN(g10764) );
AND2_X4 U_g11347 ( .A1(g6232), .A2(g213), .ZN(g11347) );
AND2_X4 U_g11420 ( .A1(g6314), .A2(g216), .ZN(g11420) );
AND2_X4 U_g11421 ( .A1(g6232), .A2(g222), .ZN(g11421) );
AND2_X4 U_g11431 ( .A1(g6369), .A2(g900), .ZN(g11431) );
AND2_X4 U_g11607 ( .A1(g5871), .A2(g8360), .ZN(g11607) );
AND2_X4 U_g11612 ( .A1(g5881), .A2(g8378), .ZN(g11612) );
AND2_X4 U_g11637 ( .A1(g5918), .A2(g8427), .ZN(g11637) );
AND2_X4 U_g11771 ( .A1(g554), .A2(g8622), .ZN(g11771) );
AND2_X4 U_g11788 ( .A1(g1240), .A2(g8632), .ZN(g11788) );
AND2_X4 U_g11805 ( .A1(g6173), .A2(g8643), .ZN(g11805) );
AND2_X4 U_g11814 ( .A1(g1934), .A2(g8651), .ZN(g11814) );
AND2_X4 U_g11816 ( .A1(g7869), .A2(g8655), .ZN(g11816) );
AND2_X4 U_g11838 ( .A1(g6205), .A2(g8659), .ZN(g11838) );
AND2_X4 U_g11847 ( .A1(g2628), .A2(g8667), .ZN(g11847) );
AND2_X4 U_g11851 ( .A1(g7849), .A2(g8670), .ZN(g11851) );
AND2_X4 U_g11880 ( .A1(g6294), .A2(g8678), .ZN(g11880) );
AND2_X4 U_g11885 ( .A1(g7834), .A2(g8684), .ZN(g11885) );
AND2_X4 U_g11922 ( .A1(g6431), .A2(g8690), .ZN(g11922) );
AND2_X4 U_g11926 ( .A1(g8169), .A2(g8696), .ZN(g11926) );
AND2_X4 U_g11966 ( .A1(g8090), .A2(g8708), .ZN(g11966) );
AND2_X4 U_g11967 ( .A1(g7967), .A2(g8711), .ZN(g11967) );
AND2_X4 U_g12012 ( .A1(g8015), .A2(g8745), .ZN(g12012) );
AND2_X4 U_g12069 ( .A1(g7964), .A2(g8763), .ZN(g12069) );
AND2_X4 U_g12070 ( .A1(g8018), .A2(g8766), .ZN(g12070) );
AND2_X4 U_g12128 ( .A1(g7916), .A2(g8785), .ZN(g12128) );
AND2_X4 U_g12129 ( .A1(g7872), .A2(g8788), .ZN(g12129) );
AND2_X4 U_g12186 ( .A1(g8093), .A2(g8805), .ZN(g12186) );
AND2_X4 U_g12273 ( .A1(g8172), .A2(g8829), .ZN(g12273) );
AND2_X4 U_g12274 ( .A1(g7900), .A2(g8832), .ZN(g12274) );
AND2_X4 U_g12307 ( .A1(g7919), .A2(g8853), .ZN(g12307) );
AND2_X4 U_g12330 ( .A1(g8246), .A2(g8879), .ZN(g12330) );
AND2_X4 U_g12331 ( .A1(g7927), .A2(g8882), .ZN(g12331) );
AND2_X4 U_g12353 ( .A1(g7852), .A2(g8915), .ZN(g12353) );
AND2_X4 U_g12376 ( .A1(g7974), .A2(g8949), .ZN(g12376) );
AND2_X4 U_g12419 ( .A1(g8028), .A2(g9006), .ZN(g12419) );
AND2_X4 U_g12429 ( .A1(g8101), .A2(g9044), .ZN(g12429) );
AND2_X4 U_g12477 ( .A1(g7822), .A2(g9128), .ZN(g12477) );
AND2_X4 U_g12494 ( .A1(g7833), .A2(g9134), .ZN(g12494) );
AND2_X4 U_g12514 ( .A1(g7848), .A2(g9140), .ZN(g12514) );
AND2_X4 U_g12531 ( .A1(g7868), .A2(g9146), .ZN(g12531) );
AND2_X4 U_g12650 ( .A1(g6149), .A2(g9290), .ZN(g12650) );
AND4_X4 U_I19937 ( .A1(g9507), .A2(g9427), .A3(g9356), .A4(g9293), .ZN(I19937) );
AND4_X4 U_I19938 ( .A1(g9232), .A2(g9187), .A3(g9161), .A4(g9150), .ZN(I19938) );
AND2_X4 U_g12876 ( .A1(I19937), .A2(I19938), .ZN(g12876) );
AND2_X4 U_g12908 ( .A1(g7899), .A2(g10004), .ZN(g12908) );
AND4_X4 U_I19971 ( .A1(g9649), .A2(g9569), .A3(g9453), .A4(g9374), .ZN(I19971) );
AND4_X4 U_I19972 ( .A1(g9310), .A2(g9248), .A3(g9203), .A4(g9174), .ZN(I19972) );
AND2_X4 U_g12916 ( .A1(I19971), .A2(I19972), .ZN(g12916) );
AND2_X4 U_g12938 ( .A1(g8179), .A2(g10096), .ZN(g12938) );
AND4_X4 U_I19996 ( .A1(g9795), .A2(g9711), .A3(g9595), .A4(g9471), .ZN(I19996) );
AND4_X4 U_I19997 ( .A1(g9391), .A2(g9326), .A3(g9264), .A4(g9216), .ZN(I19997) );
AND2_X4 U_g12945 ( .A1(I19996), .A2(I19997), .ZN(g12945) );
AND2_X4 U_g12966 ( .A1(g7926), .A2(g10189), .ZN(g12966) );
AND4_X4 U_I20021 ( .A1(g9941), .A2(g9857), .A3(g9737), .A4(g9613), .ZN(I20021) );
AND4_X4 U_I20022 ( .A1(g9488), .A2(g9407), .A3(g9342), .A4(g9277), .ZN(I20022) );
AND2_X4 U_g12974 ( .A1(I20021), .A2(I20022), .ZN(g12974) );
AND2_X4 U_g12989 ( .A1(g8254), .A2(g10273), .ZN(g12989) );
AND2_X4 U_g12990 ( .A1(g8180), .A2(g10276), .ZN(g12990) );
AND2_X4 U_g13000 ( .A1(g7973), .A2(g10357), .ZN(g13000) );
AND2_X4 U_g13004 ( .A1(g10186), .A2(g8317), .ZN(g13004) );
AND2_X4 U_g13009 ( .A1(g3995), .A2(g10416), .ZN(g13009) );
AND2_X4 U_g13010 ( .A1(g8255), .A2(g10419), .ZN(g13010) );
AND2_X4 U_g13023 ( .A1(g8027), .A2(g10482), .ZN(g13023) );
AND2_X4 U_g13031 ( .A1(g7879), .A2(g10542), .ZN(g13031) );
AND2_X4 U_g13032 ( .A1(g3996), .A2(g10545), .ZN(g13032) );
AND2_X4 U_g13042 ( .A1(g8100), .A2(g10601), .ZN(g13042) );
AND3_X4 U_I20100 ( .A1(g10186), .A2(g3018), .A3(g3028), .ZN(I20100) );
AND3_X4 U_g13055 ( .A1(g7471), .A2(g7570), .A3(I20100), .ZN(g13055) );
AND2_X4 U_g13056 ( .A1(g4092), .A2(g10646), .ZN(g13056) );
AND4_X4 U_I20131 ( .A1(g8313), .A2(g7542), .A3(g2888), .A4(g7566), .ZN(I20131) );
AND4_X4 U_I20132 ( .A1(g2892), .A2(g2903), .A3(g7595), .A4(g2908), .ZN(I20132) );
AND2_X4 U_g13082 ( .A1(I20131), .A2(I20132), .ZN(g13082) );
AND4_X4 U_g13110 ( .A1(g10693), .A2(g2883), .A3(g7562), .A4(g10711), .ZN(g13110) );
AND2_X4 U_g13247 ( .A1(g298), .A2(g11032), .ZN(g13247) );
AND2_X4 U_g13266 ( .A1(g5628), .A2(g11088), .ZN(g13266) );
AND2_X4 U_g13270 ( .A1(g985), .A2(g11102), .ZN(g13270) );
AND2_X4 U_g13289 ( .A1(g5647), .A2(g11141), .ZN(g13289) );
AND2_X4 U_g13291 ( .A1(g5656), .A2(g11154), .ZN(g13291) );
AND2_X4 U_g13295 ( .A1(g1679), .A2(g11170), .ZN(g13295) );
AND2_X4 U_g13316 ( .A1(g5675), .A2(g11210), .ZN(g13316) );
AND2_X4 U_g13320 ( .A1(g5685), .A2(g11225), .ZN(g13320) );
AND2_X4 U_g13322 ( .A1(g5694), .A2(g11240), .ZN(g13322) );
AND2_X4 U_g13326 ( .A1(g2373), .A2(g11256), .ZN(g13326) );
AND2_X4 U_g13335 ( .A1(g5708), .A2(g11278), .ZN(g13335) );
AND2_X4 U_g13340 ( .A1(g5727), .A2(g11294), .ZN(g13340) );
AND2_X4 U_g13343 ( .A1(g5737), .A2(g11309), .ZN(g13343) );
AND2_X4 U_g13345 ( .A1(g5746), .A2(g11324), .ZN(g13345) );
AND2_X4 U_g13355 ( .A1(g5756), .A2(g11355), .ZN(g13355) );
AND2_X4 U_g13360 ( .A1(g5766), .A2(g11373), .ZN(g13360) );
AND2_X4 U_g13365 ( .A1(g5785), .A2(g11389), .ZN(g13365) );
AND2_X4 U_g13368 ( .A1(g5795), .A2(g11404), .ZN(g13368) );
AND2_X4 U_g13385 ( .A1(g5815), .A2(g11441), .ZN(g13385) );
AND2_X4 U_g13390 ( .A1(g5825), .A2(g11459), .ZN(g13390) );
AND2_X4 U_g13395 ( .A1(g5844), .A2(g11475), .ZN(g13395) );
AND2_X4 U_g13477 ( .A1(g6016), .A2(g12191), .ZN(g13477) );
AND2_X4 U_g13479 ( .A1(g6017), .A2(g12196), .ZN(g13479) );
AND2_X4 U_g13480 ( .A1(g6018), .A2(g12197), .ZN(g13480) );
AND2_X4 U_g13481 ( .A1(g5864), .A2(g11603), .ZN(g13481) );
AND2_X4 U_g13483 ( .A1(g6020), .A2(g12209), .ZN(g13483) );
AND2_X4 U_g13484 ( .A1(g6021), .A2(g12210), .ZN(g13484) );
AND2_X4 U_g13485 ( .A1(g6022), .A2(g12211), .ZN(g13485) );
AND2_X4 U_g13486 ( .A1(g6023), .A2(g12212), .ZN(g13486) );
AND2_X4 U_g13487 ( .A1(g5874), .A2(g11608), .ZN(g13487) );
AND2_X4 U_g13488 ( .A1(g6025), .A2(g12218), .ZN(g13488) );
AND2_X4 U_g13489 ( .A1(g6026), .A2(g12219), .ZN(g13489) );
AND2_X4 U_g13490 ( .A1(g6027), .A2(g12220), .ZN(g13490) );
AND2_X4 U_g13491 ( .A1(g6028), .A2(g12221), .ZN(g13491) );
AND2_X4 U_g13492 ( .A1(g2371), .A2(g12222), .ZN(g13492) );
AND2_X4 U_g13493 ( .A1(g5887), .A2(g11613), .ZN(g13493) );
AND2_X4 U_g13496 ( .A1(g6032), .A2(g12246), .ZN(g13496) );
AND2_X4 U_g13498 ( .A1(g6033), .A2(g12251), .ZN(g13498) );
AND2_X4 U_g13499 ( .A1(g6034), .A2(g12252), .ZN(g13499) );
AND2_X4 U_g13500 ( .A1(g5911), .A2(g11633), .ZN(g13500) );
AND2_X4 U_g13502 ( .A1(g6036), .A2(g12264), .ZN(g13502) );
AND2_X4 U_g13503 ( .A1(g6037), .A2(g12265), .ZN(g13503) );
AND2_X4 U_g13504 ( .A1(g6038), .A2(g12266), .ZN(g13504) );
AND2_X4 U_g13505 ( .A1(g6039), .A2(g12267), .ZN(g13505) );
AND2_X4 U_g13506 ( .A1(g5921), .A2(g11638), .ZN(g13506) );
AND2_X4 U_g13513 ( .A1(g6043), .A2(g12289), .ZN(g13513) );
AND2_X4 U_g13515 ( .A1(g6044), .A2(g12294), .ZN(g13515) );
AND2_X4 U_g13516 ( .A1(g6045), .A2(g12295), .ZN(g13516) );
AND2_X4 U_g13517 ( .A1(g5950), .A2(g11656), .ZN(g13517) );
AND2_X4 U_g13527 ( .A1(g6047), .A2(g12325), .ZN(g13527) );
AND2_X4 U_g13609 ( .A1(g6141), .A2(g12456), .ZN(g13609) );
AND2_X4 U_g13619 ( .A1(g6162), .A2(g12466), .ZN(g13619) );
AND2_X4 U_g13623 ( .A1(g5428), .A2(g12472), .ZN(g13623) );
AND2_X4 U_g13625 ( .A1(g6173), .A2(g12476), .ZN(g13625) );
AND2_X4 U_g13631 ( .A1(g6189), .A2(g12481), .ZN(g13631) );
AND2_X4 U_g13634 ( .A1(g12776), .A2(g8617), .ZN(g13634) );
AND2_X4 U_g13636 ( .A1(g6205), .A2(g12493), .ZN(g13636) );
AND2_X4 U_g13642 ( .A1(g6221), .A2(g12498), .ZN(g13642) );
AND2_X4 U_g13643 ( .A1(g5431), .A2(g12502), .ZN(g13643) );
AND2_X4 U_g13645 ( .A1(g6281), .A2(g12504), .ZN(g13645) );
AND2_X4 U_g13646 ( .A1(g7772), .A2(g12505), .ZN(g13646) );
AND2_X4 U_g13648 ( .A1(g6294), .A2(g12513), .ZN(g13648) );
AND2_X4 U_g13654 ( .A1(g8093), .A2(g11791), .ZN(g13654) );
AND2_X4 U_g13655 ( .A1(g7540), .A2(g12518), .ZN(g13655) );
AND2_X4 U_g13656 ( .A1(g12776), .A2(g8640), .ZN(g13656) );
AND2_X4 U_g13671 ( .A1(g6418), .A2(g12521), .ZN(g13671) );
AND2_X4 U_g13672 ( .A1(g7788), .A2(g12522), .ZN(g13672) );
AND2_X4 U_g13674 ( .A1(g6431), .A2(g12530), .ZN(g13674) );
AND2_X4 U_g13675 ( .A1(g7561), .A2(g12532), .ZN(g13675) );
AND2_X4 U_g13676 ( .A1(g5434), .A2(g12533), .ZN(g13676) );
AND2_X4 U_g13701 ( .A1(g6623), .A2(g12536), .ZN(g13701) );
AND2_X4 U_g13702 ( .A1(g7802), .A2(g12537), .ZN(g13702) );
AND2_X4 U_g13703 ( .A1(g8018), .A2(g11848), .ZN(g13703) );
AND2_X4 U_g13704 ( .A1(g7581), .A2(g12542), .ZN(g13704) );
AND2_X4 U_g13705 ( .A1(g12776), .A2(g8673), .ZN(g13705) );
AND2_X4 U_g13738 ( .A1(g6887), .A2(g12545), .ZN(g13738) );
AND2_X4 U_g13739 ( .A1(g7815), .A2(g12546), .ZN(g13739) );
AND2_X4 U_g13740 ( .A1(g6636), .A2(g12547), .ZN(g13740) );
AND2_X4 U_g13755 ( .A1(g7347), .A2(g12551), .ZN(g13755) );
AND2_X4 U_g13787 ( .A1(g7967), .A2(g11923), .ZN(g13787) );
AND2_X4 U_g13788 ( .A1(g6897), .A2(g12553), .ZN(g13788) );
AND2_X4 U_g13789 ( .A1(g7140), .A2(g12554), .ZN(g13789) );
AND2_X4 U_g13790 ( .A1(g7475), .A2(g12558), .ZN(g13790) );
AND2_X4 U_g13796 ( .A1(g7477), .A2(g12559), .ZN(g13796) );
AND2_X4 U_g13815 ( .A1(g7139), .A2(g12560), .ZN(g13815) );
AND2_X4 U_g13816 ( .A1(g7530), .A2(g12596), .ZN(g13816) );
AND2_X4 U_g13818 ( .A1(g7531), .A2(g12597), .ZN(g13818) );
AND2_X4 U_g13824 ( .A1(g7533), .A2(g12598), .ZN(g13824) );
AND2_X4 U_g13833 ( .A1(g7919), .A2(g12009), .ZN(g13833) );
AND2_X4 U_g13834 ( .A1(g7336), .A2(g12599), .ZN(g13834) );
AND2_X4 U_g13835 ( .A1(g7461), .A2(g12600), .ZN(g13835) );
AND2_X4 U_g13837 ( .A1(g7556), .A2(g12642), .ZN(g13837) );
AND2_X4 U_g13839 ( .A1(g7557), .A2(g12643), .ZN(g13839) );
AND2_X4 U_g13845 ( .A1(g7559), .A2(g12644), .ZN(g13845) );
AND2_X4 U_g13846 ( .A1(g7460), .A2(g12645), .ZN(g13846) );
AND2_X4 U_g13847 ( .A1(g7521), .A2(g12646), .ZN(g13847) );
AND2_X4 U_g13851 ( .A1(g7579), .A2(g12688), .ZN(g13851) );
AND2_X4 U_g13853 ( .A1(g7580), .A2(g12689), .ZN(g13853) );
AND2_X4 U_g13854 ( .A1(g5349), .A2(g12690), .ZN(g13854) );
AND2_X4 U_g13855 ( .A1(g7541), .A2(g12691), .ZN(g13855) );
AND2_X4 U_g13860 ( .A1(g7593), .A2(g12742), .ZN(g13860) );
AND2_X4 U_g13862 ( .A1(g5366), .A2(g12743), .ZN(g13862) );
AND2_X4 U_g13865 ( .A1(g548), .A2(g12748), .ZN(g13865) );
AND2_X4 U_g13870 ( .A1(g7582), .A2(g12768), .ZN(g13870) );
AND2_X4 U_g13871 ( .A1(g7898), .A2(g12775), .ZN(g13871) );
AND2_X4 U_g13878 ( .A1(g7610), .A2(g12782), .ZN(g13878) );
AND2_X4 U_g13880 ( .A1(g1234), .A2(g12790), .ZN(g13880) );
AND2_X4 U_g13884 ( .A1(g7594), .A2(g12807), .ZN(g13884) );
AND2_X4 U_g13892 ( .A1(g7616), .A2(g12815), .ZN(g13892) );
AND2_X4 U_g13900 ( .A1(g7619), .A2(g12821), .ZN(g13900) );
AND2_X4 U_g13902 ( .A1(g1928), .A2(g12829), .ZN(g13902) );
AND2_X4 U_g13904 ( .A1(g7337), .A2(g12843), .ZN(g13904) );
AND2_X4 U_g13905 ( .A1(g7925), .A2(g12847), .ZN(g13905) );
AND2_X4 U_g13913 ( .A1(g7623), .A2(g12850), .ZN(g13913) );
AND2_X4 U_g13914 ( .A1(g7626), .A2(g12851), .ZN(g13914) );
AND2_X4 U_g13933 ( .A1(g7632), .A2(g12853), .ZN(g13933) );
AND2_X4 U_g13941 ( .A1(g7635), .A2(g12859), .ZN(g13941) );
AND2_X4 U_g13943 ( .A1(g2622), .A2(g12867), .ZN(g13943) );
AND2_X4 U_g13944 ( .A1(g7141), .A2(g12874), .ZN(g13944) );
AND2_X4 U_g13952 ( .A1(g7643), .A2(g12881), .ZN(g13952) );
AND2_X4 U_g13953 ( .A1(g7646), .A2(g12882), .ZN(g13953) );
AND2_X4 U_g13969 ( .A1(g7652), .A2(g12891), .ZN(g13969) );
AND2_X4 U_g13970 ( .A1(g7655), .A2(g12892), .ZN(g13970) );
AND2_X4 U_g13989 ( .A1(g7661), .A2(g12894), .ZN(g13989) );
AND2_X4 U_g13997 ( .A1(g7664), .A2(g12900), .ZN(g13997) );
AND2_X4 U_g13998 ( .A1(g7972), .A2(g12907), .ZN(g13998) );
AND2_X4 U_g14006 ( .A1(g7670), .A2(g12914), .ZN(g14006) );
AND2_X4 U_g14007 ( .A1(g7673), .A2(g12915), .ZN(g14007) );
AND2_X4 U_g14022 ( .A1(g7679), .A2(g12921), .ZN(g14022) );
AND2_X4 U_g14023 ( .A1(g7682), .A2(g12922), .ZN(g14023) );
AND2_X4 U_g14039 ( .A1(g7688), .A2(g12931), .ZN(g14039) );
AND2_X4 U_g14040 ( .A1(g7691), .A2(g12932), .ZN(g14040) );
AND2_X4 U_g14059 ( .A1(g7697), .A2(g12934), .ZN(g14059) );
AND2_X4 U_g14067 ( .A1(g7703), .A2(g12940), .ZN(g14067) );
AND2_X4 U_g14097 ( .A1(g7706), .A2(g12943), .ZN(g14097) );
AND2_X4 U_g14098 ( .A1(g7709), .A2(g12944), .ZN(g14098) );
AND2_X4 U_g14113 ( .A1(g7715), .A2(g12950), .ZN(g14113) );
AND2_X4 U_g14114 ( .A1(g7718), .A2(g12951), .ZN(g14114) );
AND2_X4 U_g14130 ( .A1(g7724), .A2(g12960), .ZN(g14130) );
AND2_X4 U_g14131 ( .A1(g7727), .A2(g12961), .ZN(g14131) );
AND2_X4 U_g14143 ( .A1(g8026), .A2(g12965), .ZN(g14143) );
AND2_X4 U_g14182 ( .A1(g7733), .A2(g12969), .ZN(g14182) );
AND2_X4 U_g14212 ( .A1(g7736), .A2(g12972), .ZN(g14212) );
AND2_X4 U_g14213 ( .A1(g7739), .A2(g12973), .ZN(g14213) );
AND2_X4 U_g14228 ( .A1(g7745), .A2(g12979), .ZN(g14228) );
AND2_X4 U_g14229 ( .A1(g7748), .A2(g12980), .ZN(g14229) );
AND2_X4 U_g14297 ( .A1(g7757), .A2(g12993), .ZN(g14297) );
AND2_X4 U_g14327 ( .A1(g7760), .A2(g12996), .ZN(g14327) );
AND2_X4 U_g14328 ( .A1(g7763), .A2(g12997), .ZN(g14328) );
AND2_X4 U_g14336 ( .A1(g8099), .A2(g12998), .ZN(g14336) );
AND2_X4 U_g14419 ( .A1(g7779), .A2(g13003), .ZN(g14419) );
AND2_X4 U_g14690 ( .A1(g7841), .A2(g13101), .ZN(g14690) );
AND2_X4 U_g14724 ( .A1(g7861), .A2(g13117), .ZN(g14724) );
AND2_X4 U_g14752 ( .A1(g7891), .A2(g13130), .ZN(g14752) );
AND2_X4 U_g14767 ( .A1(g13245), .A2(g10765), .ZN(g14767) );
AND2_X4 U_g14773 ( .A1(g7915), .A2(g13141), .ZN(g14773) );
AND2_X4 U_g14884 ( .A1(g8169), .A2(g12548), .ZN(g14884) );
AND2_X4 U_g14894 ( .A1(g3940), .A2(g13148), .ZN(g14894) );
AND2_X4 U_g14956 ( .A1(g11059), .A2(g13151), .ZN(g14956) );
AND2_X4 U_g14957 ( .A1(g4015), .A2(g13152), .ZN(g14957) );
AND2_X4 U_g14958 ( .A1(g4016), .A2(g13153), .ZN(g14958) );
AND2_X4 U_g14975 ( .A1(g4047), .A2(g13154), .ZN(g14975) );
AND2_X4 U_g15020 ( .A1(g8090), .A2(g12561), .ZN(g15020) );
AND2_X4 U_g15030 ( .A1(g4110), .A2(g13158), .ZN(g15030) );
AND2_X4 U_g15031 ( .A1(g4111), .A2(g13159), .ZN(g15031) );
AND2_X4 U_g15046 ( .A1(g4142), .A2(g13161), .ZN(g15046) );
AND2_X4 U_g15047 ( .A1(g4143), .A2(g13162), .ZN(g15047) );
AND2_X4 U_g15064 ( .A1(g4174), .A2(g13163), .ZN(g15064) );
AND2_X4 U_g15093 ( .A1(g7869), .A2(g12601), .ZN(g15093) );
AND2_X4 U_g15094 ( .A1(g7872), .A2(g12604), .ZN(g15094) );
AND2_X4 U_g15104 ( .A1(g4220), .A2(g13167), .ZN(g15104) );
AND2_X4 U_g15105 ( .A1(g4224), .A2(g13168), .ZN(g15105) );
AND2_X4 U_g15126 ( .A1(g4249), .A2(g13169), .ZN(g15126) );
AND2_X4 U_g15127 ( .A1(g4250), .A2(g13170), .ZN(g15127) );
AND2_X4 U_g15142 ( .A1(g4281), .A2(g13172), .ZN(g15142) );
AND2_X4 U_g15143 ( .A1(g4282), .A2(g13173), .ZN(g15143) );
AND2_X4 U_g15160 ( .A1(g4313), .A2(g13174), .ZN(g15160) );
AND2_X4 U_g15171 ( .A1(g8015), .A2(g12647), .ZN(g15171) );
AND2_X4 U_g15172 ( .A1(g4346), .A2(g13176), .ZN(g15172) );
AND2_X4 U_g15173 ( .A1(g4347), .A2(g13177), .ZN(g15173) );
AND2_X4 U_g15178 ( .A1(g640), .A2(g12651), .ZN(g15178) );
AND2_X4 U_g15196 ( .A1(g4375), .A2(g13178), .ZN(g15196) );
AND2_X4 U_g15197 ( .A1(g4379), .A2(g13179), .ZN(g15197) );
AND2_X4 U_g15218 ( .A1(g4404), .A2(g13180), .ZN(g15218) );
AND2_X4 U_g15219 ( .A1(g4405), .A2(g13181), .ZN(g15219) );
AND2_X4 U_g15234 ( .A1(g4436), .A2(g13183), .ZN(g15234) );
AND2_X4 U_g15235 ( .A1(g4437), .A2(g13184), .ZN(g15235) );
AND2_X4 U_g15243 ( .A1(g7849), .A2(g12692), .ZN(g15243) );
AND2_X4 U_g15244 ( .A1(g7852), .A2(g12695), .ZN(g15244) );
AND2_X4 U_g15245 ( .A1(g4474), .A2(g13185), .ZN(g15245) );
AND2_X4 U_g15246 ( .A1(g4475), .A2(g13186), .ZN(g15246) );
AND2_X4 U_g15247 ( .A1(g4479), .A2(g13187), .ZN(g15247) );
AND2_X4 U_g15257 ( .A1(g4357), .A2(g12702), .ZN(g15257) );
AND2_X4 U_g15258 ( .A1(g4515), .A2(g13188), .ZN(g15258) );
AND2_X4 U_g15259 ( .A1(g4516), .A2(g13189), .ZN(g15259) );
AND2_X4 U_g15264 ( .A1(g1326), .A2(g12705), .ZN(g15264) );
AND2_X4 U_g15282 ( .A1(g4544), .A2(g13190), .ZN(g15282) );
AND2_X4 U_g15283 ( .A1(g4548), .A2(g13191), .ZN(g15283) );
AND2_X4 U_g15304 ( .A1(g4573), .A2(g13192), .ZN(g15304) );
AND2_X4 U_g15305 ( .A1(g4574), .A2(g13193), .ZN(g15305) );
AND2_X4 U_g15320 ( .A1(g7964), .A2(g12744), .ZN(g15320) );
AND2_X4 U_g15321 ( .A1(g4601), .A2(g13195), .ZN(g15321) );
AND2_X4 U_g15324 ( .A1(g4609), .A2(g13196), .ZN(g15324) );
AND2_X4 U_g15325 ( .A1(g4610), .A2(g13197), .ZN(g15325) );
AND2_X4 U_g15335 ( .A1(g4489), .A2(g12749), .ZN(g15335) );
AND2_X4 U_g15336 ( .A1(g4492), .A2(g12752), .ZN(g15336) );
AND2_X4 U_g15337 ( .A1(g4650), .A2(g13198), .ZN(g15337) );
AND2_X4 U_g15338 ( .A1(g4651), .A2(g13199), .ZN(g15338) );
AND2_X4 U_g15339 ( .A1(g4655), .A2(g13200), .ZN(g15339) );
AND2_X4 U_g15349 ( .A1(g4526), .A2(g12759), .ZN(g15349) );
AND2_X4 U_g15350 ( .A1(g4691), .A2(g13201), .ZN(g15350) );
AND2_X4 U_g15351 ( .A1(g4692), .A2(g13202), .ZN(g15351) );
AND2_X4 U_g15356 ( .A1(g2020), .A2(g12762), .ZN(g15356) );
AND2_X4 U_g15374 ( .A1(g4720), .A2(g13203), .ZN(g15374) );
AND2_X4 U_g15375 ( .A1(g4724), .A2(g13204), .ZN(g15375) );
AND2_X4 U_g15388 ( .A1(g7834), .A2(g12769), .ZN(g15388) );
AND2_X4 U_g15389 ( .A1(g8246), .A2(g12772), .ZN(g15389) );
AND2_X4 U_g15391 ( .A1(g4752), .A2(g13205), .ZN(g15391) );
AND2_X4 U_g15392 ( .A1(g4753), .A2(g13206), .ZN(g15392) );
AND2_X4 U_g15402 ( .A1(g4620), .A2(g12783), .ZN(g15402) );
AND2_X4 U_g15403 ( .A1(g4623), .A2(g12786), .ZN(g15403) );
AND2_X4 U_g15407 ( .A1(g4778), .A2(g13207), .ZN(g15407) );
AND2_X4 U_g15410 ( .A1(g4786), .A2(g13208), .ZN(g15410) );
AND2_X4 U_g15411 ( .A1(g4787), .A2(g13209), .ZN(g15411) );
AND2_X4 U_g15421 ( .A1(g4665), .A2(g12791), .ZN(g15421) );
AND2_X4 U_g15422 ( .A1(g4668), .A2(g12794), .ZN(g15422) );
AND2_X4 U_g15423 ( .A1(g4827), .A2(g13210), .ZN(g15423) );
AND2_X4 U_g15424 ( .A1(g4828), .A2(g13211), .ZN(g15424) );
AND2_X4 U_g15425 ( .A1(g4832), .A2(g13212), .ZN(g15425) );
AND2_X4 U_g15435 ( .A1(g4702), .A2(g12801), .ZN(g15435) );
AND2_X4 U_g15436 ( .A1(g4868), .A2(g13213), .ZN(g15436) );
AND2_X4 U_g15437 ( .A1(g4869), .A2(g13214), .ZN(g15437) );
AND2_X4 U_g15442 ( .A1(g2714), .A2(g12804), .ZN(g15442) );
AND2_X4 U_g15452 ( .A1(g7916), .A2(g12808), .ZN(g15452) );
AND2_X4 U_g15453 ( .A1(g6898), .A2(g12811), .ZN(g15453) );
AND2_X4 U_g15459 ( .A1(g4897), .A2(g13218), .ZN(g15459) );
AND2_X4 U_g15460 ( .A1(g4898), .A2(g13219), .ZN(g15460) );
AND2_X4 U_g15470 ( .A1(g4763), .A2(g12816), .ZN(g15470) );
AND2_X4 U_g15475 ( .A1(g4928), .A2(g13220), .ZN(g15475) );
AND2_X4 U_g15476 ( .A1(g4929), .A2(g13221), .ZN(g15476) );
AND2_X4 U_g15486 ( .A1(g4797), .A2(g12822), .ZN(g15486) );
AND2_X4 U_g15487 ( .A1(g4800), .A2(g12825), .ZN(g15487) );
AND2_X4 U_g15491 ( .A1(g4954), .A2(g13222), .ZN(g15491) );
AND2_X4 U_g15494 ( .A1(g4962), .A2(g13223), .ZN(g15494) );
AND2_X4 U_g15495 ( .A1(g4963), .A2(g13224), .ZN(g15495) );
AND2_X4 U_g15505 ( .A1(g4842), .A2(g12830), .ZN(g15505) );
AND2_X4 U_g15506 ( .A1(g4845), .A2(g12833), .ZN(g15506) );
AND2_X4 U_g15507 ( .A1(g5003), .A2(g13225), .ZN(g15507) );
AND2_X4 U_g15508 ( .A1(g5004), .A2(g13226), .ZN(g15508) );
AND2_X4 U_g15509 ( .A1(g5008), .A2(g13227), .ZN(g15509) );
AND2_X4 U_g15519 ( .A1(g4879), .A2(g12840), .ZN(g15519) );
AND2_X4 U_g15520 ( .A1(g8172), .A2(g12844), .ZN(g15520) );
AND2_X4 U_g15526 ( .A1(g5033), .A2(g13232), .ZN(g15526) );
AND2_X4 U_g15527 ( .A1(g5034), .A2(g13233), .ZN(g15527) );
AND2_X4 U_g15545 ( .A1(g5056), .A2(g13237), .ZN(g15545) );
AND2_X4 U_g15546 ( .A1(g5057), .A2(g13238), .ZN(g15546) );
AND2_X4 U_g15556 ( .A1(g4939), .A2(g12854), .ZN(g15556) );
AND2_X4 U_g15561 ( .A1(g5087), .A2(g13239), .ZN(g15561) );
AND2_X4 U_g15562 ( .A1(g5088), .A2(g13240), .ZN(g15562) );
AND2_X4 U_g15572 ( .A1(g4973), .A2(g12860), .ZN(g15572) );
AND2_X4 U_g15573 ( .A1(g4976), .A2(g12863), .ZN(g15573) );
AND2_X4 U_g15577 ( .A1(g5113), .A2(g13241), .ZN(g15577) );
AND2_X4 U_g15580 ( .A1(g5121), .A2(g13242), .ZN(g15580) );
AND2_X4 U_g15581 ( .A1(g5122), .A2(g13243), .ZN(g15581) );
AND2_X4 U_g15591 ( .A1(g5018), .A2(g12868), .ZN(g15591) );
AND2_X4 U_g15592 ( .A1(g5021), .A2(g12871), .ZN(g15592) );
AND2_X4 U_g15593 ( .A1(g7897), .A2(g13244), .ZN(g15593) );
AND2_X4 U_g15594 ( .A1(g5148), .A2(g13249), .ZN(g15594) );
AND2_X4 U_g15595 ( .A1(g5149), .A2(g13250), .ZN(g15595) );
AND2_X4 U_g15604 ( .A1(g5162), .A2(g13255), .ZN(g15604) );
AND2_X4 U_g15605 ( .A1(g5163), .A2(g13256), .ZN(g15605) );
AND2_X4 U_g15623 ( .A1(g5185), .A2(g13260), .ZN(g15623) );
AND2_X4 U_g15624 ( .A1(g5186), .A2(g13261), .ZN(g15624) );
AND2_X4 U_g15634 ( .A1(g5098), .A2(g12895), .ZN(g15634) );
AND2_X4 U_g15639 ( .A1(g5216), .A2(g13262), .ZN(g15639) );
AND2_X4 U_g15640 ( .A1(g5217), .A2(g13263), .ZN(g15640) );
AND2_X4 U_g15650 ( .A1(g5132), .A2(g12901), .ZN(g15650) );
AND2_X4 U_g15651 ( .A1(g5135), .A2(g12904), .ZN(g15651) );
AND2_X4 U_g15658 ( .A1(g8177), .A2(g13264), .ZN(g15658) );
AND2_X4 U_g15666 ( .A1(g5233), .A2(g13268), .ZN(g15666) );
AND2_X4 U_g15670 ( .A1(g5241), .A2(g13272), .ZN(g15670) );
AND2_X4 U_g15671 ( .A1(g5242), .A2(g13273), .ZN(g15671) );
AND2_X4 U_g15680 ( .A1(g5255), .A2(g13278), .ZN(g15680) );
AND2_X4 U_g15681 ( .A1(g5256), .A2(g13279), .ZN(g15681) );
AND2_X4 U_g15699 ( .A1(g5278), .A2(g13283), .ZN(g15699) );
AND2_X4 U_g15700 ( .A1(g5279), .A2(g13284), .ZN(g15700) );
AND2_X4 U_g15710 ( .A1(g5227), .A2(g12935), .ZN(g15710) );
AND2_X4 U_g15717 ( .A1(g7924), .A2(g13285), .ZN(g15717) );
AND2_X4 U_g15725 ( .A1(g5296), .A2(g13293), .ZN(g15725) );
AND2_X4 U_g15729 ( .A1(g5304), .A2(g13297), .ZN(g15729) );
AND2_X4 U_g15730 ( .A1(g5305), .A2(g13298), .ZN(g15730) );
AND2_X4 U_g15739 ( .A1(g5318), .A2(g13303), .ZN(g15739) );
AND2_X4 U_g15740 ( .A1(g5319), .A2(g13304), .ZN(g15740) );
AND2_X4 U_g15753 ( .A1(g7542), .A2(g12962), .ZN(g15753) );
AND2_X4 U_g15754 ( .A1(g7837), .A2(g13308), .ZN(g15754) );
AND2_X4 U_g15755 ( .A1(g8178), .A2(g13309), .ZN(g15755) );
AND2_X4 U_g15765 ( .A1(g5333), .A2(g13324), .ZN(g15765) );
AND2_X4 U_g15769 ( .A1(g5341), .A2(g13328), .ZN(g15769) );
AND2_X4 U_g15770 ( .A1(g5342), .A2(g13329), .ZN(g15770) );
AND3_X4 U_I22028 ( .A1(g13004), .A2(g3018), .A3(g7549), .ZN(I22028) );
AND3_X4 U_g15780 ( .A1(g7471), .A2(g3032), .A3(I22028), .ZN(g15780) );
AND2_X4 U_g15781 ( .A1(g7971), .A2(g13330), .ZN(g15781) );
AND2_X4 U_g15793 ( .A1(g5361), .A2(g13347), .ZN(g15793) );
AND2_X4 U_g15801 ( .A1(g7856), .A2(g13351), .ZN(g15801) );
AND2_X4 U_g15802 ( .A1(g8253), .A2(g13352), .ZN(g15802) );
AND2_X4 U_g15817 ( .A1(g8025), .A2(g13373), .ZN(g15817) );
AND2_X4 U_g15828 ( .A1(g7877), .A2(g13398), .ZN(g15828) );
AND2_X4 U_g15829 ( .A1(g7857), .A2(g13400), .ZN(g15829) );
AND2_X4 U_g15840 ( .A1(g8098), .A2(g11620), .ZN(g15840) );
AND2_X4 U_g15852 ( .A1(g7878), .A2(g11642), .ZN(g15852) );
AND3_X4 U_I22136 ( .A1(g13082), .A2(g2912), .A3(g7522), .ZN(I22136) );
AND3_X4 U_g15902 ( .A1(g7607), .A2(g2920), .A3(I22136), .ZN(g15902) );
AND2_X4 U_g15998 ( .A1(g5469), .A2(g11732), .ZN(g15998) );
AND2_X4 U_g16003 ( .A1(g12013), .A2(g10826), .ZN(g16003) );
AND2_X4 U_g16004 ( .A1(g5587), .A2(g11734), .ZN(g16004) );
AND2_X4 U_g16008 ( .A1(g5504), .A2(g11735), .ZN(g16008) );
AND2_X4 U_g16009 ( .A1(g12071), .A2(g10843), .ZN(g16009) );
AND2_X4 U_g16010 ( .A1(g7639), .A2(g11736), .ZN(g16010) );
AND2_X4 U_g16015 ( .A1(g12013), .A2(g10859), .ZN(g16015) );
AND2_X4 U_g16016 ( .A1(g5601), .A2(g11740), .ZN(g16016) );
AND2_X4 U_g16017 ( .A1(g12130), .A2(g10862), .ZN(g16017) );
AND2_X4 U_g16018 ( .A1(g6149), .A2(g11741), .ZN(g16018) );
AND2_X4 U_g16019 ( .A1(g5507), .A2(g11742), .ZN(g16019) );
AND2_X4 U_g16028 ( .A1(g5543), .A2(g11745), .ZN(g16028) );
AND2_X4 U_g16029 ( .A1(g12071), .A2(g10877), .ZN(g16029) );
AND2_X4 U_g16030 ( .A1(g7667), .A2(g11746), .ZN(g16030) );
AND2_X4 U_g16031 ( .A1(g6227), .A2(g11747), .ZN(g16031) );
AND2_X4 U_g16032 ( .A1(g12187), .A2(g10883), .ZN(g16032) );
AND2_X4 U_g16033 ( .A1(g5546), .A2(g11748), .ZN(g16033) );
AND2_X4 U_g16045 ( .A1(g12013), .A2(g10892), .ZN(g16045) );
AND2_X4 U_g16046 ( .A1(g5618), .A2(g11761), .ZN(g16046) );
AND2_X4 U_g16047 ( .A1(g12130), .A2(g10895), .ZN(g16047) );
AND2_X4 U_g16048 ( .A1(g6170), .A2(g11762), .ZN(g16048) );
AND2_X4 U_g16049 ( .A1(g6638), .A2(g11763), .ZN(g16049) );
AND2_X4 U_g16050 ( .A1(g5590), .A2(g11764), .ZN(g16050) );
AND2_X4 U_g16051 ( .A1(g12235), .A2(g10901), .ZN(g16051) );
AND2_X4 U_g16052 ( .A1(g5591), .A2(g11765), .ZN(g16052) );
AND2_X4 U_g16053 ( .A1(g297), .A2(g11770), .ZN(g16053) );
AND2_X4 U_g16066 ( .A1(g12071), .A2(g10912), .ZN(g16066) );
AND2_X4 U_g16067 ( .A1(g7700), .A2(g11774), .ZN(g16067) );
AND2_X4 U_g16068 ( .A1(g6310), .A2(g11775), .ZN(g16068) );
AND2_X4 U_g16069 ( .A1(g5346), .A2(g11776), .ZN(g16069) );
AND2_X4 U_g16070 ( .A1(g12187), .A2(g10921), .ZN(g16070) );
AND2_X4 U_g16071 ( .A1(g5604), .A2(g11777), .ZN(g16071) );
AND2_X4 U_g16072 ( .A1(g12275), .A2(g10924), .ZN(g16072) );
AND2_X4 U_g16073 ( .A1(g5605), .A2(g11778), .ZN(g16073) );
AND2_X4 U_g16074 ( .A1(g5646), .A2(g11782), .ZN(g16074) );
AND2_X4 U_g16081 ( .A1(g3304), .A2(g11783), .ZN(g16081) );
AND2_X4 U_g16089 ( .A1(g984), .A2(g11787), .ZN(g16089) );
AND2_X4 U_g16100 ( .A1(g12130), .A2(g10937), .ZN(g16100) );
AND2_X4 U_g16101 ( .A1(g6197), .A2(g11794), .ZN(g16101) );
AND2_X4 U_g16102 ( .A1(g6905), .A2(g11795), .ZN(g16102) );
AND2_X4 U_g16103 ( .A1(g5621), .A2(g11796), .ZN(g16103) );
AND2_X4 U_g16104 ( .A1(g12235), .A2(g10946), .ZN(g16104) );
AND2_X4 U_g16105 ( .A1(g5622), .A2(g11797), .ZN(g16105) );
AND2_X4 U_g16106 ( .A1(g12308), .A2(g10949), .ZN(g16106) );
AND2_X4 U_g16107 ( .A1(g5666), .A2(g11801), .ZN(g16107) );
AND2_X4 U_g16108 ( .A1(g5667), .A2(g11802), .ZN(g16108) );
AND2_X4 U_g16109 ( .A1(g8277), .A2(g11803), .ZN(g16109) );
AND2_X4 U_g16110 ( .A1(g516), .A2(g11804), .ZN(g16110) );
AND2_X4 U_g16111 ( .A1(g5551), .A2(g13215), .ZN(g16111) );
AND2_X4 U_g16112 ( .A1(g5684), .A2(g11808), .ZN(g16112) );
AND2_X4 U_g16119 ( .A1(g3460), .A2(g11809), .ZN(g16119) );
AND2_X4 U_g16127 ( .A1(g1678), .A2(g11813), .ZN(g16127) );
AND2_X4 U_g16133 ( .A1(g6444), .A2(g11817), .ZN(g16133) );
AND2_X4 U_g16134 ( .A1(g5363), .A2(g11818), .ZN(g16134) );
AND2_X4 U_g16135 ( .A1(g12187), .A2(g10980), .ZN(g16135) );
AND2_X4 U_g16136 ( .A1(g5640), .A2(g11819), .ZN(g16136) );
AND2_X4 U_g16137 ( .A1(g12275), .A2(g10983), .ZN(g16137) );
AND2_X4 U_g16138 ( .A1(g5641), .A2(g11820), .ZN(g16138) );
AND2_X4 U_g16139 ( .A1(g5704), .A2(g11824), .ZN(g16139) );
AND2_X4 U_g16140 ( .A1(g5705), .A2(g11825), .ZN(g16140) );
AND2_X4 U_g16141 ( .A1(g5706), .A2(g11826), .ZN(g16141) );
AND2_X4 U_g16152 ( .A1(g517), .A2(g11829), .ZN(g16152) );
AND2_X4 U_g16153 ( .A1(g5592), .A2(g13229), .ZN(g16153) );
AND2_X4 U_g16158 ( .A1(g5718), .A2(g11834), .ZN(g16158) );
AND2_X4 U_g16159 ( .A1(g5719), .A2(g11835), .ZN(g16159) );
AND2_X4 U_g16160 ( .A1(g8286), .A2(g11836), .ZN(g16160) );
AND2_X4 U_g16161 ( .A1(g1202), .A2(g11837), .ZN(g16161) );
AND2_X4 U_g16162 ( .A1(g5597), .A2(g13234), .ZN(g16162) );
AND2_X4 U_g16163 ( .A1(g5736), .A2(g11841), .ZN(g16163) );
AND2_X4 U_g16170 ( .A1(g3616), .A2(g11842), .ZN(g16170) );
AND2_X4 U_g16178 ( .A1(g2372), .A2(g11846), .ZN(g16178) );
AND2_X4 U_g16182 ( .A1(g7149), .A2(g11852), .ZN(g16182) );
AND2_X4 U_g16183 ( .A1(g12235), .A2(g11014), .ZN(g16183) );
AND2_X4 U_g16184 ( .A1(g5663), .A2(g11853), .ZN(g16184) );
AND2_X4 U_g16185 ( .A1(g12308), .A2(g11017), .ZN(g16185) );
AND2_X4 U_g16186 ( .A1(g5753), .A2(g11856), .ZN(g16186) );
AND2_X4 U_g16187 ( .A1(g5754), .A2(g11857), .ZN(g16187) );
AND2_X4 U_g16188 ( .A1(g5755), .A2(g11858), .ZN(g16188) );
AND2_X4 U_g16197 ( .A1(g518), .A2(g11862), .ZN(g16197) );
AND2_X4 U_g16198 ( .A1(g5762), .A2(g11866), .ZN(g16198) );
AND2_X4 U_g16199 ( .A1(g5763), .A2(g11867), .ZN(g16199) );
AND2_X4 U_g16200 ( .A1(g5764), .A2(g11868), .ZN(g16200) );
AND2_X4 U_g16211 ( .A1(g1203), .A2(g11871), .ZN(g16211) );
AND2_X4 U_g16212 ( .A1(g5609), .A2(g13252), .ZN(g16212) );
AND2_X4 U_g16217 ( .A1(g5776), .A2(g11876), .ZN(g16217) );
AND2_X4 U_g16218 ( .A1(g5777), .A2(g11877), .ZN(g16218) );
AND2_X4 U_g16219 ( .A1(g8295), .A2(g11878), .ZN(g16219) );
AND2_X4 U_g16220 ( .A1(g1896), .A2(g11879), .ZN(g16220) );
AND2_X4 U_g16221 ( .A1(g5614), .A2(g13257), .ZN(g16221) );
AND2_X4 U_g16222 ( .A1(g5794), .A2(g11883), .ZN(g16222) );
AND2_X4 U_g16229 ( .A1(g3772), .A2(g11884), .ZN(g16229) );
AND2_X4 U_g16237 ( .A1(g5379), .A2(g11886), .ZN(g16237) );
AND2_X4 U_g16238 ( .A1(g12275), .A2(g11066), .ZN(g16238) );
AND2_X4 U_g16239 ( .A1(g5700), .A2(g11887), .ZN(g16239) );
AND2_X4 U_g16240 ( .A1(g5804), .A2(g11891), .ZN(g16240) );
AND2_X4 U_g16241 ( .A1(g5805), .A2(g11892), .ZN(g16241) );
AND2_X4 U_g16242 ( .A1(g5806), .A2(g11893), .ZN(g16242) );
AND2_X4 U_g16250 ( .A1(g519), .A2(g11895), .ZN(g16250) );
AND2_X4 U_g16251 ( .A1(g5812), .A2(g11898), .ZN(g16251) );
AND2_X4 U_g16252 ( .A1(g5813), .A2(g11899), .ZN(g16252) );
AND2_X4 U_g16253 ( .A1(g5814), .A2(g11900), .ZN(g16253) );
AND2_X4 U_g16262 ( .A1(g1204), .A2(g11904), .ZN(g16262) );
AND2_X4 U_g16263 ( .A1(g5821), .A2(g11908), .ZN(g16263) );
AND2_X4 U_g16264 ( .A1(g5822), .A2(g11909), .ZN(g16264) );
AND2_X4 U_g16265 ( .A1(g5823), .A2(g11910), .ZN(g16265) );
AND2_X4 U_g16276 ( .A1(g1897), .A2(g11913), .ZN(g16276) );
AND2_X4 U_g16277 ( .A1(g5634), .A2(g13275), .ZN(g16277) );
AND2_X4 U_g16282 ( .A1(g5835), .A2(g11918), .ZN(g16282) );
AND2_X4 U_g16283 ( .A1(g5836), .A2(g11919), .ZN(g16283) );
AND2_X4 U_g16284 ( .A1(g8304), .A2(g11920), .ZN(g16284) );
AND2_X4 U_g16285 ( .A1(g2590), .A2(g11921), .ZN(g16285) );
AND2_X4 U_g16286 ( .A1(g5639), .A2(g13280), .ZN(g16286) );
AND2_X4 U_g16288 ( .A1(g12308), .A2(g11129), .ZN(g16288) );
AND2_X4 U_g16289 ( .A1(g5853), .A2(g11929), .ZN(g16289) );
AND2_X4 U_g16290 ( .A1(g5854), .A2(g11930), .ZN(g16290) );
AND2_X4 U_g16291 ( .A1(g5855), .A2(g11931), .ZN(g16291) );
AND2_X4 U_g16292 ( .A1(g294), .A2(g11932), .ZN(g16292) );
AND2_X4 U_g16298 ( .A1(g520), .A2(g11936), .ZN(g16298) );
AND2_X4 U_g16299 ( .A1(g5860), .A2(g11941), .ZN(g16299) );
AND2_X4 U_g16300 ( .A1(g5861), .A2(g11942), .ZN(g16300) );
AND2_X4 U_g16301 ( .A1(g5862), .A2(g11943), .ZN(g16301) );
AND2_X4 U_g16309 ( .A1(g1205), .A2(g11945), .ZN(g16309) );
AND2_X4 U_g16310 ( .A1(g5868), .A2(g11948), .ZN(g16310) );
AND2_X4 U_g16311 ( .A1(g5869), .A2(g11949), .ZN(g16311) );
AND2_X4 U_g16312 ( .A1(g5870), .A2(g11950), .ZN(g16312) );
AND2_X4 U_g16321 ( .A1(g1898), .A2(g11954), .ZN(g16321) );
AND2_X4 U_g16322 ( .A1(g5877), .A2(g11958), .ZN(g16322) );
AND2_X4 U_g16323 ( .A1(g5878), .A2(g11959), .ZN(g16323) );
AND2_X4 U_g16324 ( .A1(g5879), .A2(g11960), .ZN(g16324) );
AND2_X4 U_g16335 ( .A1(g2591), .A2(g11963), .ZN(g16335) );
AND2_X4 U_g16336 ( .A1(g5662), .A2(g13300), .ZN(g16336) );
AND2_X4 U_g16342 ( .A1(g5894), .A2(g11968), .ZN(g16342) );
AND2_X4 U_g16343 ( .A1(g5895), .A2(g11969), .ZN(g16343) );
AND2_X4 U_g16344 ( .A1(g5896), .A2(g11970), .ZN(g16344) );
AND2_X4 U_g16345 ( .A1(g5897), .A2(g11971), .ZN(g16345) );
AND2_X4 U_g16346 ( .A1(g295), .A2(g11972), .ZN(g16346) );
AND2_X4 U_g16347 ( .A1(g5900), .A2(g11982), .ZN(g16347) );
AND2_X4 U_g16348 ( .A1(g5901), .A2(g11983), .ZN(g16348) );
AND2_X4 U_g16349 ( .A1(g5902), .A2(g11984), .ZN(g16349) );
AND2_X4 U_g16350 ( .A1(g981), .A2(g11985), .ZN(g16350) );
AND2_X4 U_g16356 ( .A1(g1206), .A2(g11989), .ZN(g16356) );
AND2_X4 U_g16357 ( .A1(g5907), .A2(g11994), .ZN(g16357) );
AND2_X4 U_g16358 ( .A1(g5908), .A2(g11995), .ZN(g16358) );
AND2_X4 U_g16359 ( .A1(g5909), .A2(g11996), .ZN(g16359) );
AND2_X4 U_g16367 ( .A1(g1899), .A2(g11998), .ZN(g16367) );
AND2_X4 U_g16368 ( .A1(g5915), .A2(g12001), .ZN(g16368) );
AND2_X4 U_g16369 ( .A1(g5916), .A2(g12002), .ZN(g16369) );
AND2_X4 U_g16370 ( .A1(g5917), .A2(g12003), .ZN(g16370) );
AND2_X4 U_g16379 ( .A1(g2592), .A2(g12007), .ZN(g16379) );
AND2_X4 U_g16380 ( .A1(g5925), .A2(g12020), .ZN(g16380) );
AND2_X4 U_g16381 ( .A1(g5926), .A2(g12021), .ZN(g16381) );
AND2_X4 U_g16382 ( .A1(g5927), .A2(g12022), .ZN(g16382) );
AND2_X4 U_g16383 ( .A1(g5928), .A2(g12023), .ZN(g16383) );
AND2_X4 U_g16384 ( .A1(g296), .A2(g12024), .ZN(g16384) );
AND2_X4 U_g16385 ( .A1(g5714), .A2(g13336), .ZN(g16385) );
AND2_X4 U_g16386 ( .A1(g5933), .A2(g12037), .ZN(g16386) );
AND2_X4 U_g16387 ( .A1(g5934), .A2(g12038), .ZN(g16387) );
AND2_X4 U_g16388 ( .A1(g5935), .A2(g12039), .ZN(g16388) );
AND2_X4 U_g16389 ( .A1(g5936), .A2(g12040), .ZN(g16389) );
AND2_X4 U_g16390 ( .A1(g982), .A2(g12041), .ZN(g16390) );
AND2_X4 U_g16391 ( .A1(g5939), .A2(g12051), .ZN(g16391) );
AND2_X4 U_g16392 ( .A1(g5940), .A2(g12052), .ZN(g16392) );
AND2_X4 U_g16393 ( .A1(g5941), .A2(g12053), .ZN(g16393) );
AND2_X4 U_g16394 ( .A1(g1675), .A2(g12054), .ZN(g16394) );
AND2_X4 U_g16400 ( .A1(g1900), .A2(g12058), .ZN(g16400) );
AND2_X4 U_g16401 ( .A1(g5946), .A2(g12063), .ZN(g16401) );
AND2_X4 U_g16402 ( .A1(g5947), .A2(g12064), .ZN(g16402) );
AND2_X4 U_g16403 ( .A1(g5948), .A2(g12065), .ZN(g16403) );
AND2_X4 U_g16411 ( .A1(g2593), .A2(g12067), .ZN(g16411) );
AND2_X4 U_g16413 ( .A1(g5954), .A2(g12075), .ZN(g16413) );
AND2_X4 U_g16414 ( .A1(g5955), .A2(g12076), .ZN(g16414) );
AND2_X4 U_g16415 ( .A1(g5956), .A2(g12077), .ZN(g16415) );
AND2_X4 U_g16416 ( .A1(g5957), .A2(g12078), .ZN(g16416) );
AND2_X4 U_g16417 ( .A1(g5759), .A2(g13356), .ZN(g16417) );
AND2_X4 U_g16418 ( .A1(g5959), .A2(g12084), .ZN(g16418) );
AND2_X4 U_g16419 ( .A1(g5960), .A2(g12085), .ZN(g16419) );
AND2_X4 U_g16420 ( .A1(g5961), .A2(g12086), .ZN(g16420) );
AND2_X4 U_g16421 ( .A1(g5962), .A2(g12087), .ZN(g16421) );
AND2_X4 U_g16422 ( .A1(g983), .A2(g12088), .ZN(g16422) );
AND2_X4 U_g16423 ( .A1(g5772), .A2(g13361), .ZN(g16423) );
AND2_X4 U_g16424 ( .A1(g5967), .A2(g12101), .ZN(g16424) );
AND2_X4 U_g16425 ( .A1(g5968), .A2(g12102), .ZN(g16425) );
AND2_X4 U_g16426 ( .A1(g5969), .A2(g12103), .ZN(g16426) );
AND2_X4 U_g16427 ( .A1(g5970), .A2(g12104), .ZN(g16427) );
AND2_X4 U_g16428 ( .A1(g1676), .A2(g12105), .ZN(g16428) );
AND2_X4 U_g16429 ( .A1(g5973), .A2(g12115), .ZN(g16429) );
AND2_X4 U_g16430 ( .A1(g5974), .A2(g12116), .ZN(g16430) );
AND2_X4 U_g16431 ( .A1(g5975), .A2(g12117), .ZN(g16431) );
AND2_X4 U_g16432 ( .A1(g2369), .A2(g12118), .ZN(g16432) );
AND2_X4 U_g16438 ( .A1(g2594), .A2(g12122), .ZN(g16438) );
AND2_X4 U_g16443 ( .A1(g5980), .A2(g12134), .ZN(g16443) );
AND2_X4 U_g16444 ( .A1(g5981), .A2(g12135), .ZN(g16444) );
AND2_X4 U_g16445 ( .A1(g5808), .A2(g13381), .ZN(g16445) );
AND2_X4 U_g16447 ( .A1(g5983), .A2(g12147), .ZN(g16447) );
AND2_X4 U_g16448 ( .A1(g5984), .A2(g12148), .ZN(g16448) );
AND2_X4 U_g16449 ( .A1(g5985), .A2(g12149), .ZN(g16449) );
AND2_X4 U_g16450 ( .A1(g5986), .A2(g12150), .ZN(g16450) );
AND2_X4 U_g16451 ( .A1(g5818), .A2(g13386), .ZN(g16451) );
AND2_X4 U_g16452 ( .A1(g5988), .A2(g12156), .ZN(g16452) );
AND2_X4 U_g16453 ( .A1(g5989), .A2(g12157), .ZN(g16453) );
AND2_X4 U_g16454 ( .A1(g5990), .A2(g12158), .ZN(g16454) );
AND2_X4 U_g16455 ( .A1(g5991), .A2(g12159), .ZN(g16455) );
AND2_X4 U_g16456 ( .A1(g1677), .A2(g12160), .ZN(g16456) );
AND2_X4 U_g16457 ( .A1(g5831), .A2(g13391), .ZN(g16457) );
AND2_X4 U_g16458 ( .A1(g5996), .A2(g12173), .ZN(g16458) );
AND2_X4 U_g16459 ( .A1(g5997), .A2(g12174), .ZN(g16459) );
AND2_X4 U_g16460 ( .A1(g5998), .A2(g12175), .ZN(g16460) );
AND2_X4 U_g16461 ( .A1(g5999), .A2(g12176), .ZN(g16461) );
AND2_X4 U_g16462 ( .A1(g2370), .A2(g12177), .ZN(g16462) );
AND4_X4 U_g16505 ( .A1(g14776), .A2(g14797), .A3(g16142), .A4(g16243), .ZN(g16505) );
AND4_X4 U_g16513 ( .A1(g15065), .A2(g13724), .A3(g13764), .A4(g13797), .ZN(g16513) );
AND4_X4 U_g16527 ( .A1(g14811), .A2(g14849), .A3(g16201), .A4(g16302), .ZN(g16527) );
AND4_X4 U_g16535 ( .A1(g15161), .A2(g13774), .A3(g13805), .A4(g13825), .ZN(g16535) );
AND4_X4 U_g16558 ( .A1(g14863), .A2(g14922), .A3(g16266), .A4(g16360), .ZN(g16558) );
AND4_X4 U_g16590 ( .A1(g14936), .A2(g15003), .A3(g16325), .A4(g16404), .ZN(g16590) );
AND2_X4 U_g16607 ( .A1(g15022), .A2(g15096), .ZN(g16607) );
AND2_X4 U_g16625 ( .A1(g15118), .A2(g15188), .ZN(g16625) );
AND2_X4 U_g16639 ( .A1(g15210), .A2(g15274), .ZN(g16639) );
AND2_X4 U_g16650 ( .A1(g15296), .A2(g15366), .ZN(g16650) );
AND2_X4 U_g16850 ( .A1(g6226), .A2(g14764), .ZN(g16850) );
AND2_X4 U_g16855 ( .A1(g15722), .A2(g8646), .ZN(g16855) );
AND2_X4 U_g16856 ( .A1(g6443), .A2(g14794), .ZN(g16856) );
AND2_X4 U_g16859 ( .A1(g15762), .A2(g8662), .ZN(g16859) );
AND2_X4 U_g16864 ( .A1(g15790), .A2(g8681), .ZN(g16864) );
AND2_X4 U_g16865 ( .A1(g6896), .A2(g14881), .ZN(g16865) );
AND2_X4 U_g16879 ( .A1(g15813), .A2(g8693), .ZN(g16879) );
AND2_X4 U_g16894 ( .A1(g7156), .A2(g14959), .ZN(g16894) );
AND2_X4 U_g16907 ( .A1(g7335), .A2(g15017), .ZN(g16907) );
AND2_X4 U_g16908 ( .A1(g7838), .A2(g15032), .ZN(g16908) );
AND2_X4 U_g16909 ( .A1(g6908), .A2(g15033), .ZN(g16909) );
AND2_X4 U_g16923 ( .A1(g7352), .A2(g15048), .ZN(g16923) );
AND2_X4 U_g16938 ( .A1(g7858), .A2(g15128), .ZN(g16938) );
AND2_X4 U_g16939 ( .A1(g7158), .A2(g15129), .ZN(g16939) );
AND2_X4 U_g16953 ( .A1(g7482), .A2(g15144), .ZN(g16953) );
AND2_X4 U_g16964 ( .A1(g7520), .A2(g15170), .ZN(g16964) );
AND2_X4 U_g16966 ( .A1(g7529), .A2(g15174), .ZN(g16966) );
AND2_X4 U_g16967 ( .A1(g7827), .A2(g15175), .ZN(g16967) );
AND2_X4 U_g16968 ( .A1(g6672), .A2(g15176), .ZN(g16968) );
AND2_X4 U_g16969 ( .A1(g7888), .A2(g15220), .ZN(g16969) );
AND2_X4 U_g16970 ( .A1(g7354), .A2(g15221), .ZN(g16970) );
AND2_X4 U_g16984 ( .A1(g7538), .A2(g15236), .ZN(g16984) );
AND2_X4 U_g16987 ( .A1(g7555), .A2(g15260), .ZN(g16987) );
AND2_X4 U_g16988 ( .A1(g7842), .A2(g15261), .ZN(g16988) );
AND2_X4 U_g16989 ( .A1(g6974), .A2(g15262), .ZN(g16989) );
AND2_X4 U_g16990 ( .A1(g7912), .A2(g15306), .ZN(g16990) );
AND2_X4 U_g16991 ( .A1(g7484), .A2(g15307), .ZN(g16991) );
AND2_X4 U_g16993 ( .A1(g7576), .A2(g15322), .ZN(g16993) );
AND2_X4 U_g16994 ( .A1(g7819), .A2(g15323), .ZN(g16994) );
AND2_X4 U_g16997 ( .A1(g7578), .A2(g15352), .ZN(g16997) );
AND2_X4 U_g16998 ( .A1(g7862), .A2(g15353), .ZN(g16998) );
AND2_X4 U_g16999 ( .A1(g7224), .A2(g15354), .ZN(g16999) );
AND3_X4 U_g17001 ( .A1(g3254), .A2(g10694), .A3(g14144), .ZN(g17001) );
AND2_X4 U_g17015 ( .A1(g7996), .A2(g15390), .ZN(g17015) );
AND2_X4 U_g17017 ( .A1(g7590), .A2(g15408), .ZN(g17017) );
AND2_X4 U_g17018 ( .A1(g7830), .A2(g15409), .ZN(g17018) );
AND2_X4 U_g17021 ( .A1(g7592), .A2(g15438), .ZN(g17021) );
AND2_X4 U_g17022 ( .A1(g7892), .A2(g15439), .ZN(g17022) );
AND2_X4 U_g17023 ( .A1(g7420), .A2(g15440), .ZN(g17023) );
AND2_X4 U_g17028 ( .A1(g7604), .A2(g15458), .ZN(g17028) );
AND3_X4 U_g17031 ( .A1(g3410), .A2(g10714), .A3(g14259), .ZN(g17031) );
AND2_X4 U_g17045 ( .A1(g8071), .A2(g15474), .ZN(g17045) );
AND2_X4 U_g17047 ( .A1(g7605), .A2(g15492), .ZN(g17047) );
AND2_X4 U_g17048 ( .A1(g7845), .A2(g15493), .ZN(g17048) );
AND2_X4 U_g17055 ( .A1(g7153), .A2(g15524), .ZN(g17055) );
AND2_X4 U_g17056 ( .A1(g7953), .A2(g15525), .ZN(g17056) );
AND2_X4 U_g17062 ( .A1(g7613), .A2(g15544), .ZN(g17062) );
AND3_X4 U_g17065 ( .A1(g3566), .A2(g10735), .A3(g14381), .ZN(g17065) );
AND2_X4 U_g17079 ( .A1(g8156), .A2(g15560), .ZN(g17079) );
AND2_X4 U_g17081 ( .A1(g7614), .A2(g15578), .ZN(g17081) );
AND2_X4 U_g17082 ( .A1(g7865), .A2(g15579), .ZN(g17082) );
AND2_X4 U_g17084 ( .A1(g7629), .A2(g13954), .ZN(g17084) );
AND2_X4 U_g17090 ( .A1(g7349), .A2(g15602), .ZN(g17090) );
AND2_X4 U_g17091 ( .A1(g8004), .A2(g15603), .ZN(g17091) );
AND2_X4 U_g17097 ( .A1(g7622), .A2(g15622), .ZN(g17097) );
AND3_X4 U_g17100 ( .A1(g3722), .A2(g10754), .A3(g14493), .ZN(g17100) );
AND2_X4 U_g17114 ( .A1(g8242), .A2(g15638), .ZN(g17114) );
AND2_X4 U_g17116 ( .A1(g7649), .A2(g14008), .ZN(g17116) );
AND2_X4 U_g17117 ( .A1(g7906), .A2(g15665), .ZN(g17117) );
AND2_X4 U_g17122 ( .A1(g7658), .A2(g14024), .ZN(g17122) );
AND2_X4 U_g17128 ( .A1(g7479), .A2(g15678), .ZN(g17128) );
AND2_X4 U_g17129 ( .A1(g8079), .A2(g15679), .ZN(g17129) );
AND2_X4 U_g17135 ( .A1(g7638), .A2(g15698), .ZN(g17135) );
AND2_X4 U_g17138 ( .A1(g7676), .A2(g14068), .ZN(g17138) );
AND2_X4 U_g17143 ( .A1(g7685), .A2(g14099), .ZN(g17143) );
AND2_X4 U_g17144 ( .A1(g7958), .A2(g15724), .ZN(g17144) );
AND2_X4 U_g17149 ( .A1(g7694), .A2(g14115), .ZN(g17149) );
AND2_X4 U_g17155 ( .A1(g7535), .A2(g15737), .ZN(g17155) );
AND2_X4 U_g17156 ( .A1(g8164), .A2(g15738), .ZN(g17156) );
AND2_X4 U_g17161 ( .A1(g7712), .A2(g14183), .ZN(g17161) );
AND2_X4 U_g17166 ( .A1(g7721), .A2(g14214), .ZN(g17166) );
AND2_X4 U_g17167 ( .A1(g8009), .A2(g15764), .ZN(g17167) );
AND2_X4 U_g17172 ( .A1(g7730), .A2(g14230), .ZN(g17172) );
AND2_X4 U_g17176 ( .A1(g7742), .A2(g14298), .ZN(g17176) );
AND2_X4 U_g17181 ( .A1(g7751), .A2(g14329), .ZN(g17181) );
AND2_X4 U_g17182 ( .A1(g8084), .A2(g15792), .ZN(g17182) );
AND2_X4 U_g17193 ( .A1(g7766), .A2(g14420), .ZN(g17193) );
AND2_X4 U_g17268 ( .A1(g8024), .A2(g15991), .ZN(g17268) );
AND2_X4 U_g17301 ( .A1(g8097), .A2(g15994), .ZN(g17301) );
AND2_X4 U_g17339 ( .A1(g8176), .A2(g15997), .ZN(g17339) );
AND2_X4 U_g17352 ( .A1(g3942), .A2(g14960), .ZN(g17352) );
AND2_X4 U_g17353 ( .A1(g3945), .A2(g14963), .ZN(g17353) );
AND2_X4 U_g17381 ( .A1(g8250), .A2(g16001), .ZN(g17381) );
AND2_X4 U_g17382 ( .A1(g8252), .A2(g16002), .ZN(g17382) );
AND2_X4 U_g17393 ( .A1(g3941), .A2(g16005), .ZN(g17393) );
AND2_X4 U_g17395 ( .A1(g6177), .A2(g15034), .ZN(g17395) );
AND2_X4 U_g17396 ( .A1(g4020), .A2(g15037), .ZN(g17396) );
AND2_X4 U_g17397 ( .A1(g4023), .A2(g15040), .ZN(g17397) );
AND2_X4 U_g17398 ( .A1(g4026), .A2(g15043), .ZN(g17398) );
AND2_X4 U_g17408 ( .A1(g4049), .A2(g15049), .ZN(g17408) );
AND2_X4 U_g17409 ( .A1(g4052), .A2(g15052), .ZN(g17409) );
AND2_X4 U_g17428 ( .A1(g3994), .A2(g16007), .ZN(g17428) );
AND2_X4 U_g17446 ( .A1(g6284), .A2(g16011), .ZN(g17446) );
AND2_X4 U_g17447 ( .A1(g4115), .A2(g15106), .ZN(g17447) );
AND2_X4 U_g17448 ( .A1(g4118), .A2(g15109), .ZN(g17448) );
AND2_X4 U_g17449 ( .A1(g4121), .A2(g15112), .ZN(g17449) );
AND2_X4 U_g17450 ( .A1(g4124), .A2(g15115), .ZN(g17450) );
AND2_X4 U_g17460 ( .A1(g4048), .A2(g16012), .ZN(g17460) );
AND2_X4 U_g17461 ( .A1(g6209), .A2(g15130), .ZN(g17461) );
AND2_X4 U_g17462 ( .A1(g4147), .A2(g15133), .ZN(g17462) );
AND2_X4 U_g17463 ( .A1(g4150), .A2(g15136), .ZN(g17463) );
AND2_X4 U_g17464 ( .A1(g4153), .A2(g15139), .ZN(g17464) );
AND2_X4 U_g17474 ( .A1(g4176), .A2(g15145), .ZN(g17474) );
AND2_X4 U_g17475 ( .A1(g4179), .A2(g15148), .ZN(g17475) );
AND2_X4 U_g17485 ( .A1(g4089), .A2(g16013), .ZN(g17485) );
AND2_X4 U_g17486 ( .A1(g4091), .A2(g16014), .ZN(g17486) );
AND2_X4 U_g17506 ( .A1(g6675), .A2(g16023), .ZN(g17506) );
AND2_X4 U_g17508 ( .A1(g4225), .A2(g15179), .ZN(g17508) );
AND2_X4 U_g17509 ( .A1(g4228), .A2(g15182), .ZN(g17509) );
AND2_X4 U_g17510 ( .A1(g4231), .A2(g15185), .ZN(g17510) );
AND2_X4 U_g17526 ( .A1(g6421), .A2(g16025), .ZN(g17526) );
AND2_X4 U_g17527 ( .A1(g4254), .A2(g15198), .ZN(g17527) );
AND2_X4 U_g17528 ( .A1(g4257), .A2(g15201), .ZN(g17528) );
AND2_X4 U_g17529 ( .A1(g4260), .A2(g15204), .ZN(g17529) );
AND2_X4 U_g17530 ( .A1(g4263), .A2(g15207), .ZN(g17530) );
AND2_X4 U_g17540 ( .A1(g4175), .A2(g16026), .ZN(g17540) );
AND2_X4 U_g17541 ( .A1(g6298), .A2(g15222), .ZN(g17541) );
AND2_X4 U_g17542 ( .A1(g4286), .A2(g15225), .ZN(g17542) );
AND2_X4 U_g17543 ( .A1(g4289), .A2(g15228), .ZN(g17543) );
AND2_X4 U_g17544 ( .A1(g4292), .A2(g15231), .ZN(g17544) );
AND2_X4 U_g17554 ( .A1(g4315), .A2(g15237), .ZN(g17554) );
AND2_X4 U_g17555 ( .A1(g4318), .A2(g15240), .ZN(g17555) );
AND2_X4 U_g17556 ( .A1(g4201), .A2(g16027), .ZN(g17556) );
AND2_X4 U_g17576 ( .A1(g4348), .A2(g15248), .ZN(g17576) );
AND2_X4 U_g17577 ( .A1(g4351), .A2(g15251), .ZN(g17577) );
AND2_X4 U_g17578 ( .A1(g4354), .A2(g15254), .ZN(g17578) );
AND2_X4 U_g17597 ( .A1(g6977), .A2(g16039), .ZN(g17597) );
AND2_X4 U_g17598 ( .A1(g4380), .A2(g15265), .ZN(g17598) );
AND2_X4 U_g17599 ( .A1(g4383), .A2(g15268), .ZN(g17599) );
AND2_X4 U_g17600 ( .A1(g4386), .A2(g15271), .ZN(g17600) );
AND2_X4 U_g17616 ( .A1(g6626), .A2(g16041), .ZN(g17616) );
AND2_X4 U_g17617 ( .A1(g4409), .A2(g15284), .ZN(g17617) );
AND2_X4 U_g17618 ( .A1(g4412), .A2(g15287), .ZN(g17618) );
AND2_X4 U_g17619 ( .A1(g4415), .A2(g15290), .ZN(g17619) );
AND2_X4 U_g17620 ( .A1(g4418), .A2(g15293), .ZN(g17620) );
AND2_X4 U_g17630 ( .A1(g4314), .A2(g16042), .ZN(g17630) );
AND2_X4 U_g17631 ( .A1(g6435), .A2(g15308), .ZN(g17631) );
AND2_X4 U_g17632 ( .A1(g4441), .A2(g15311), .ZN(g17632) );
AND2_X4 U_g17633 ( .A1(g4444), .A2(g15314), .ZN(g17633) );
AND2_X4 U_g17634 ( .A1(g4447), .A2(g15317), .ZN(g17634) );
AND2_X4 U_g17635 ( .A1(g4322), .A2(g16043), .ZN(g17635) );
AND2_X4 U_g17636 ( .A1(g4324), .A2(g16044), .ZN(g17636) );
AND2_X4 U_g17652 ( .A1(g4480), .A2(g15326), .ZN(g17652) );
AND2_X4 U_g17653 ( .A1(g4483), .A2(g15329), .ZN(g17653) );
AND2_X4 U_g17654 ( .A1(g4486), .A2(g15332), .ZN(g17654) );
AND2_X4 U_g17673 ( .A1(g4517), .A2(g15340), .ZN(g17673) );
AND2_X4 U_g17674 ( .A1(g4520), .A2(g15343), .ZN(g17674) );
AND2_X4 U_g17675 ( .A1(g4523), .A2(g15346), .ZN(g17675) );
AND2_X4 U_g17694 ( .A1(g7227), .A2(g16061), .ZN(g17694) );
AND2_X4 U_g17695 ( .A1(g4549), .A2(g15357), .ZN(g17695) );
AND2_X4 U_g17696 ( .A1(g4552), .A2(g15360), .ZN(g17696) );
AND2_X4 U_g17697 ( .A1(g4555), .A2(g15363), .ZN(g17697) );
AND2_X4 U_g17713 ( .A1(g6890), .A2(g16063), .ZN(g17713) );
AND2_X4 U_g17714 ( .A1(g4578), .A2(g15376), .ZN(g17714) );
AND2_X4 U_g17715 ( .A1(g4581), .A2(g15379), .ZN(g17715) );
AND2_X4 U_g17716 ( .A1(g4584), .A2(g15382), .ZN(g17716) );
AND2_X4 U_g17717 ( .A1(g4587), .A2(g15385), .ZN(g17717) );
AND2_X4 U_g17718 ( .A1(g4451), .A2(g16064), .ZN(g17718) );
AND2_X4 U_g17719 ( .A1(g2993), .A2(g16065), .ZN(g17719) );
AND2_X4 U_g17734 ( .A1(g4611), .A2(g15393), .ZN(g17734) );
AND2_X4 U_g17735 ( .A1(g4614), .A2(g15396), .ZN(g17735) );
AND2_X4 U_g17736 ( .A1(g4617), .A2(g15399), .ZN(g17736) );
AND2_X4 U_g17737 ( .A1(g4626), .A2(g15404), .ZN(g17737) );
AND2_X4 U_g17752 ( .A1(g4656), .A2(g15412), .ZN(g17752) );
AND2_X4 U_g17753 ( .A1(g4659), .A2(g15415), .ZN(g17753) );
AND2_X4 U_g17754 ( .A1(g4662), .A2(g15418), .ZN(g17754) );
AND2_X4 U_g17773 ( .A1(g4693), .A2(g15426), .ZN(g17773) );
AND2_X4 U_g17774 ( .A1(g4696), .A2(g15429), .ZN(g17774) );
AND2_X4 U_g17775 ( .A1(g4699), .A2(g15432), .ZN(g17775) );
AND2_X4 U_g17794 ( .A1(g7423), .A2(g16097), .ZN(g17794) );
AND2_X4 U_g17795 ( .A1(g4725), .A2(g15443), .ZN(g17795) );
AND2_X4 U_g17796 ( .A1(g4728), .A2(g15446), .ZN(g17796) );
AND2_X4 U_g17797 ( .A1(g4731), .A2(g15449), .ZN(g17797) );
AND2_X4 U_g17798 ( .A1(g4591), .A2(g16099), .ZN(g17798) );
AND2_X4 U_g17812 ( .A1(g4754), .A2(g15461), .ZN(g17812) );
AND2_X4 U_g17813 ( .A1(g4757), .A2(g15464), .ZN(g17813) );
AND2_X4 U_g17814 ( .A1(g4760), .A2(g15467), .ZN(g17814) );
AND2_X4 U_g17824 ( .A1(g4766), .A2(g15471), .ZN(g17824) );
AND2_X4 U_g17835 ( .A1(g4788), .A2(g15477), .ZN(g17835) );
AND2_X4 U_g17836 ( .A1(g4791), .A2(g15480), .ZN(g17836) );
AND2_X4 U_g17837 ( .A1(g4794), .A2(g15483), .ZN(g17837) );
AND2_X4 U_g17838 ( .A1(g4803), .A2(g15488), .ZN(g17838) );
AND2_X4 U_g17853 ( .A1(g4833), .A2(g15496), .ZN(g17853) );
AND2_X4 U_g17854 ( .A1(g4836), .A2(g15499), .ZN(g17854) );
AND2_X4 U_g17855 ( .A1(g4839), .A2(g15502), .ZN(g17855) );
AND2_X4 U_g17874 ( .A1(g4870), .A2(g15510), .ZN(g17874) );
AND2_X4 U_g17875 ( .A1(g4873), .A2(g15513), .ZN(g17875) );
AND2_X4 U_g17876 ( .A1(g4876), .A2(g15516), .ZN(g17876) );
AND2_X4 U_g17877 ( .A1(g2998), .A2(g15521), .ZN(g17877) );
AND2_X4 U_g17900 ( .A1(g4899), .A2(g15528), .ZN(g17900) );
AND2_X4 U_g17901 ( .A1(g4902), .A2(g15531), .ZN(g17901) );
AND2_X4 U_g17902 ( .A1(g4905), .A2(g15534), .ZN(g17902) );
AND2_X4 U_g17912 ( .A1(g4908), .A2(g15537), .ZN(g17912) );
AND2_X4 U_g17924 ( .A1(g4930), .A2(g15547), .ZN(g17924) );
AND2_X4 U_g17925 ( .A1(g4933), .A2(g15550), .ZN(g17925) );
AND2_X4 U_g17926 ( .A1(g4936), .A2(g15553), .ZN(g17926) );
AND2_X4 U_g17936 ( .A1(g4942), .A2(g15557), .ZN(g17936) );
AND2_X4 U_g17947 ( .A1(g4964), .A2(g15563), .ZN(g17947) );
AND2_X4 U_g17948 ( .A1(g4967), .A2(g15566), .ZN(g17948) );
AND2_X4 U_g17949 ( .A1(g4970), .A2(g15569), .ZN(g17949) );
AND2_X4 U_g17950 ( .A1(g4979), .A2(g15574), .ZN(g17950) );
AND2_X4 U_g17965 ( .A1(g5009), .A2(g15582), .ZN(g17965) );
AND2_X4 U_g17966 ( .A1(g5012), .A2(g15585), .ZN(g17966) );
AND2_X4 U_g17967 ( .A1(g5015), .A2(g15588), .ZN(g17967) );
AND2_X4 U_g17989 ( .A1(g5035), .A2(g15596), .ZN(g17989) );
AND2_X4 U_g17990 ( .A1(g5038), .A2(g15599), .ZN(g17990) );
AND2_X4 U_g18011 ( .A1(g5058), .A2(g15606), .ZN(g18011) );
AND2_X4 U_g18012 ( .A1(g5061), .A2(g15609), .ZN(g18012) );
AND2_X4 U_g18013 ( .A1(g5064), .A2(g15612), .ZN(g18013) );
AND2_X4 U_g18023 ( .A1(g5067), .A2(g15615), .ZN(g18023) );
AND2_X4 U_g18035 ( .A1(g5089), .A2(g15625), .ZN(g18035) );
AND2_X4 U_g18036 ( .A1(g5092), .A2(g15628), .ZN(g18036) );
AND2_X4 U_g18037 ( .A1(g5095), .A2(g15631), .ZN(g18037) );
AND2_X4 U_g18047 ( .A1(g5101), .A2(g15635), .ZN(g18047) );
AND2_X4 U_g18058 ( .A1(g5123), .A2(g15641), .ZN(g18058) );
AND2_X4 U_g18059 ( .A1(g5126), .A2(g15644), .ZN(g18059) );
AND2_X4 U_g18060 ( .A1(g5129), .A2(g15647), .ZN(g18060) );
AND2_X4 U_g18061 ( .A1(g5138), .A2(g15652), .ZN(g18061) );
AND2_X4 U_g18062 ( .A1(g7462), .A2(g15655), .ZN(g18062) );
AND2_X4 U_g18088 ( .A1(g5150), .A2(g15667), .ZN(g18088) );
AND2_X4 U_g18106 ( .A1(g5164), .A2(g15672), .ZN(g18106) );
AND2_X4 U_g18107 ( .A1(g5167), .A2(g15675), .ZN(g18107) );
AND2_X4 U_g18128 ( .A1(g5187), .A2(g15682), .ZN(g18128) );
AND2_X4 U_g18129 ( .A1(g5190), .A2(g15685), .ZN(g18129) );
AND2_X4 U_g18130 ( .A1(g5193), .A2(g15688), .ZN(g18130) );
AND2_X4 U_g18140 ( .A1(g5196), .A2(g15691), .ZN(g18140) );
AND2_X4 U_g18152 ( .A1(g5218), .A2(g15701), .ZN(g18152) );
AND2_X4 U_g18153 ( .A1(g5221), .A2(g15704), .ZN(g18153) );
AND2_X4 U_g18154 ( .A1(g5224), .A2(g15707), .ZN(g18154) );
AND2_X4 U_g18164 ( .A1(g5230), .A2(g15711), .ZN(g18164) );
AND2_X4 U_g18165 ( .A1(g2883), .A2(g16287), .ZN(g18165) );
AND2_X4 U_g18169 ( .A1(g7527), .A2(g15714), .ZN(g18169) );
AND2_X4 U_g18204 ( .A1(g5243), .A2(g15726), .ZN(g18204) );
AND2_X4 U_g18222 ( .A1(g5257), .A2(g15731), .ZN(g18222) );
AND2_X4 U_g18223 ( .A1(g5260), .A2(g15734), .ZN(g18223) );
AND2_X4 U_g18244 ( .A1(g5280), .A2(g15741), .ZN(g18244) );
AND2_X4 U_g18245 ( .A1(g5283), .A2(g15744), .ZN(g18245) );
AND2_X4 U_g18246 ( .A1(g5286), .A2(g15747), .ZN(g18246) );
AND2_X4 U_g18256 ( .A1(g5289), .A2(g15750), .ZN(g18256) );
AND2_X4 U_g18311 ( .A1(g5306), .A2(g15766), .ZN(g18311) );
AND2_X4 U_g18329 ( .A1(g5320), .A2(g15771), .ZN(g18329) );
AND2_X4 U_g18330 ( .A1(g5323), .A2(g15774), .ZN(g18330) );
AND2_X4 U_g18333 ( .A1(g2888), .A2(g15777), .ZN(g18333) );
AND2_X4 U_g18404 ( .A1(g5343), .A2(g15794), .ZN(g18404) );
AND3_X4 U_I24619 ( .A1(g14776), .A2(g14837), .A3(g16142), .ZN(I24619) );
AND3_X4 U_g18547 ( .A1(g13677), .A2(g13750), .A3(I24619), .ZN(g18547) );
AND3_X4 U_I24689 ( .A1(g14811), .A2(g14910), .A3(g16201), .ZN(I24689) );
AND3_X4 U_g18597 ( .A1(g13714), .A2(g13791), .A3(I24689), .ZN(g18597) );
AND3_X4 U_I24738 ( .A1(g14863), .A2(g14991), .A3(g16266), .ZN(I24738) );
AND3_X4 U_g18629 ( .A1(g13764), .A2(g13819), .A3(I24738), .ZN(g18629) );
AND3_X4 U_I24758 ( .A1(g14936), .A2(g15080), .A3(g16325), .ZN(I24758) );
AND3_X4 U_g18638 ( .A1(g13805), .A2(g13840), .A3(I24758), .ZN(g18638) );
AND4_X4 U_g18645 ( .A1(g14776), .A2(g14895), .A3(g16142), .A4(g13750), .ZN(g18645) );
AND3_X4 U_g18647 ( .A1(g14895), .A2(g16142), .A3(g16243), .ZN(g18647) );
AND4_X4 U_g18648 ( .A1(g14811), .A2(g14976), .A3(g16201), .A4(g13791), .ZN(g18648) );
AND4_X4 U_g18649 ( .A1(g14776), .A2(g14837), .A3(g13657), .A4(g16189), .ZN(g18649) );
AND3_X4 U_g18650 ( .A1(g14976), .A2(g16201), .A3(g16302), .ZN(g18650) );
AND4_X4 U_g18651 ( .A1(g14863), .A2(g15065), .A3(g16266), .A4(g13819), .ZN(g18651) );
AND4_X4 U_g18652 ( .A1(g14797), .A2(g13657), .A3(g13677), .A4(g16243), .ZN(g18652) );
AND4_X4 U_g18653 ( .A1(g14811), .A2(g14910), .A3(g13687), .A4(g16254), .ZN(g18653) );
AND3_X4 U_g18654 ( .A1(g15065), .A2(g16266), .A3(g16360), .ZN(g18654) );
AND4_X4 U_g18655 ( .A1(g14936), .A2(g15161), .A3(g16325), .A4(g13840), .ZN(g18655) );
AND4_X4 U_g18665 ( .A1(g14776), .A2(g14837), .A3(g16189), .A4(g13706), .ZN(g18665) );
AND4_X4 U_g18666 ( .A1(g14849), .A2(g13687), .A3(g13714), .A4(g16302), .ZN(g18666) );
AND4_X4 U_g18667 ( .A1(g14863), .A2(g14991), .A3(g13724), .A4(g16313), .ZN(g18667) );
AND3_X4 U_g18668 ( .A1(g15161), .A2(g16325), .A3(g16404), .ZN(g18668) );
AND4_X4 U_g18688 ( .A1(g14811), .A2(g14910), .A3(g16254), .A4(g13756), .ZN(g18688) );
AND4_X4 U_g18689 ( .A1(g14922), .A2(g13724), .A3(g13764), .A4(g16360), .ZN(g18689) );
AND4_X4 U_g18690 ( .A1(g14936), .A2(g15080), .A3(g13774), .A4(g16371), .ZN(g18690) );
AND4_X4 U_g18717 ( .A1(g14863), .A2(g14991), .A3(g16313), .A4(g13797), .ZN(g18717) );
AND4_X4 U_g18718 ( .A1(g15003), .A2(g13774), .A3(g13805), .A4(g16404), .ZN(g18718) );
AND4_X4 U_g18753 ( .A1(g14936), .A2(g15080), .A3(g16371), .A4(g13825), .ZN(g18753) );
AND2_X4 U_g18982 ( .A1(g13519), .A2(g16154), .ZN(g18982) );
AND2_X4 U_g18990 ( .A1(g13530), .A2(g16213), .ZN(g18990) );
AND4_X4 U_g18994 ( .A1(g14895), .A2(g13657), .A3(g13677), .A4(g13706), .ZN(g18994) );
AND2_X4 U_g18997 ( .A1(g13541), .A2(g16278), .ZN(g18997) );
AND4_X4 U_g19007 ( .A1(g14976), .A2(g13687), .A3(g13714), .A4(g13756), .ZN(g19007) );
AND2_X4 U_g19010 ( .A1(g13552), .A2(g16337), .ZN(g19010) );
AND4_X4 U_g19063 ( .A1(g18679), .A2(g14910), .A3(g13687), .A4(g16254), .ZN(g19063) );
AND4_X4 U_g19079 ( .A1(g14797), .A2(g18692), .A3(g16142), .A4(g16189), .ZN(g19079) );
AND4_X4 U_g19080 ( .A1(g18708), .A2(g14991), .A3(g13724), .A4(g16313), .ZN(g19080) );
AND2_X4 U_g19087 ( .A1(g17215), .A2(g16540), .ZN(g19087) );
AND4_X4 U_g19088 ( .A1(g18656), .A2(g14797), .A3(g16189), .A4(g13706), .ZN(g19088) );
AND4_X4 U_g19089 ( .A1(g14849), .A2(g18728), .A3(g16201), .A4(g16254), .ZN(g19089) );
AND4_X4 U_g19090 ( .A1(g18744), .A2(g15080), .A3(g13774), .A4(g16371), .ZN(g19090) );
AND4_X4 U_g19092 ( .A1(g14776), .A2(g18670), .A3(g18692), .A4(g16293), .ZN(g19092) );
AND2_X4 U_g19093 ( .A1(g17218), .A2(g16572), .ZN(g19093) );
AND4_X4 U_g19094 ( .A1(g18679), .A2(g14849), .A3(g16254), .A4(g13756), .ZN(g19094) );
AND4_X4 U_g19095 ( .A1(g14922), .A2(g18765), .A3(g16266), .A4(g16313), .ZN(g19095) );
AND3_X4 U_I25280 ( .A1(g18656), .A2(g18670), .A3(g18720), .ZN(I25280) );
AND3_X4 U_g19097 ( .A1(g13657), .A2(g16243), .A3(I25280), .ZN(g19097) );
AND4_X4 U_g19099 ( .A1(g14811), .A2(g18699), .A3(g18728), .A4(g16351), .ZN(g19099) );
AND2_X4 U_g19100 ( .A1(g17220), .A2(g16596), .ZN(g19100) );
AND4_X4 U_g19101 ( .A1(g18708), .A2(g14922), .A3(g16313), .A4(g13797), .ZN(g19101) );
AND4_X4 U_g19102 ( .A1(g15003), .A2(g18796), .A3(g16325), .A4(g16371), .ZN(g19102) );
AND3_X4 U_I25291 ( .A1(g18679), .A2(g18699), .A3(g18758), .ZN(I25291) );
AND3_X4 U_g19104 ( .A1(g13687), .A2(g16302), .A3(I25291), .ZN(g19104) );
AND4_X4 U_g19106 ( .A1(g14863), .A2(g18735), .A3(g18765), .A4(g16395), .ZN(g19106) );
AND2_X4 U_g19107 ( .A1(g17223), .A2(g16616), .ZN(g19107) );
AND4_X4 U_g19108 ( .A1(g18744), .A2(g15003), .A3(g16371), .A4(g13825), .ZN(g19108) );
AND3_X4 U_I25300 ( .A1(g18708), .A2(g18735), .A3(g18789), .ZN(I25300) );
AND3_X4 U_g19109 ( .A1(g13724), .A2(g16360), .A3(I25300), .ZN(g19109) );
AND4_X4 U_g19111 ( .A1(g14936), .A2(g18772), .A3(g18796), .A4(g16433), .ZN(g19111) );
AND2_X4 U_g19112 ( .A1(g14657), .A2(g16633), .ZN(g19112) );
AND3_X4 U_I25311 ( .A1(g18744), .A2(g18772), .A3(g18815), .ZN(I25311) );
AND3_X4 U_g19116 ( .A1(g13774), .A2(g16404), .A3(I25311), .ZN(g19116) );
AND2_X4 U_g19117 ( .A1(g14691), .A2(g16644), .ZN(g19117) );
AND2_X4 U_g19124 ( .A1(g14725), .A2(g16656), .ZN(g19124) );
AND2_X4 U_g19131 ( .A1(g14753), .A2(g16673), .ZN(g19131) );
AND2_X4 U_g19142 ( .A1(g17159), .A2(g16719), .ZN(g19142) );
AND2_X4 U_g19143 ( .A1(g17174), .A2(g16761), .ZN(g19143) );
AND2_X4 U_g19146 ( .A1(g17191), .A2(g16788), .ZN(g19146) );
AND2_X4 U_g19148 ( .A1(g17202), .A2(g16817), .ZN(g19148) );
AND2_X4 U_g19150 ( .A1(g17189), .A2(g8602), .ZN(g19150) );
AND2_X4 U_g19155 ( .A1(g17200), .A2(g8614), .ZN(g19155) );
AND2_X4 U_g19161 ( .A1(g17207), .A2(g8627), .ZN(g19161) );
AND2_X4 U_g19166 ( .A1(g17212), .A2(g8637), .ZN(g19166) );
AND2_X4 U_g19228 ( .A1(g16662), .A2(g12125), .ZN(g19228) );
AND2_X4 U_g19236 ( .A1(g16935), .A2(g8802), .ZN(g19236) );
AND3_X4 U_g19241 ( .A1(g16867), .A2(g14158), .A3(g14071), .ZN(g19241) );
AND2_X4 U_g19248 ( .A1(g16662), .A2(g8817), .ZN(g19248) );
AND2_X4 U_g19252 ( .A1(g18725), .A2(g9527), .ZN(g19252) );
AND3_X4 U_g19254 ( .A1(g16895), .A2(g14273), .A3(g14186), .ZN(g19254) );
AND2_X4 U_g19260 ( .A1(g16749), .A2(g3124), .ZN(g19260) );
AND3_X4 U_g19267 ( .A1(g16924), .A2(g14395), .A3(g14301), .ZN(g19267) );
AND3_X4 U_g19282 ( .A1(g16954), .A2(g14507), .A3(g14423), .ZN(g19282) );
AND2_X4 U_g19284 ( .A1(g18063), .A2(g3111), .ZN(g19284) );
AND2_X4 U_g19285 ( .A1(g16749), .A2(g7642), .ZN(g19285) );
AND2_X4 U_g19289 ( .A1(g17029), .A2(g8580), .ZN(g19289) );
AND3_X4 U_g19303 ( .A1(g16867), .A2(g16543), .A3(g14071), .ZN(g19303) );
AND2_X4 U_g19307 ( .A1(g17063), .A2(g8587), .ZN(g19307) );
AND2_X4 U_g19316 ( .A1(g18063), .A2(g3110), .ZN(g19316) );
AND2_X4 U_g19317 ( .A1(g16749), .A2(g3126), .ZN(g19317) );
AND3_X4 U_g19320 ( .A1(g16867), .A2(g16515), .A3(g14158), .ZN(g19320) );
AND3_X4 U_g19324 ( .A1(g16895), .A2(g16575), .A3(g14186), .ZN(g19324) );
AND2_X4 U_g19328 ( .A1(g17098), .A2(g8594), .ZN(g19328) );
AND3_X4 U_g19347 ( .A1(g16895), .A2(g16546), .A3(g14273), .ZN(g19347) );
AND3_X4 U_g19351 ( .A1(g16924), .A2(g16599), .A3(g14301), .ZN(g19351) );
AND2_X4 U_g19355 ( .A1(g17136), .A2(g8605), .ZN(g19355) );
AND2_X4 U_g19356 ( .A1(g18063), .A2(g3112), .ZN(g19356) );
AND3_X4 U_g19381 ( .A1(g16924), .A2(g16578), .A3(g14395), .ZN(g19381) );
AND3_X4 U_g19385 ( .A1(g16954), .A2(g16619), .A3(g14423), .ZN(g19385) );
AND3_X4 U_g19413 ( .A1(g16954), .A2(g16602), .A3(g14507), .ZN(g19413) );
AND3_X4 U_g19449 ( .A1(g16884), .A2(g14797), .A3(g14776), .ZN(g19449) );
AND3_X4 U_g19476 ( .A1(g16913), .A2(g14849), .A3(g14811), .ZN(g19476) );
AND3_X4 U_g19499 ( .A1(g16943), .A2(g14922), .A3(g14863), .ZN(g19499) );
AND3_X4 U_g19520 ( .A1(g16974), .A2(g15003), .A3(g14936), .ZN(g19520) );
AND3_X4 U_g19531 ( .A1(g16884), .A2(g16722), .A3(g14776), .ZN(g19531) );
AND3_X4 U_g19540 ( .A1(g16884), .A2(g16697), .A3(g14797), .ZN(g19540) );
AND3_X4 U_g19541 ( .A1(g16913), .A2(g16764), .A3(g14811), .ZN(g19541) );
AND3_X4 U_g19544 ( .A1(g16913), .A2(g16728), .A3(g14849), .ZN(g19544) );
AND3_X4 U_g19545 ( .A1(g16943), .A2(g16791), .A3(g14863), .ZN(g19545) );
AND3_X4 U_g19547 ( .A1(g16943), .A2(g16770), .A3(g14922), .ZN(g19547) );
AND3_X4 U_g19548 ( .A1(g16974), .A2(g16820), .A3(g14936), .ZN(g19548) );
AND2_X4 U_g19549 ( .A1(g7950), .A2(g17230), .ZN(g19549) );
AND3_X4 U_g19551 ( .A1(g16974), .A2(g16797), .A3(g15003), .ZN(g19551) );
AND2_X4 U_g19552 ( .A1(g16829), .A2(g6048), .ZN(g19552) );
AND2_X4 U_g19553 ( .A1(g7990), .A2(g17237), .ZN(g19553) );
AND2_X4 U_g19554 ( .A1(g7993), .A2(g17240), .ZN(g19554) );
AND2_X4 U_g19555 ( .A1(g8001), .A2(g17243), .ZN(g19555) );
AND2_X4 U_g19557 ( .A1(g8053), .A2(g17249), .ZN(g19557) );
AND2_X4 U_g19558 ( .A1(g8056), .A2(g17252), .ZN(g19558) );
AND2_X4 U_g19559 ( .A1(g8059), .A2(g17255), .ZN(g19559) );
AND2_X4 U_g19560 ( .A1(g8065), .A2(g17259), .ZN(g19560) );
AND2_X4 U_g19561 ( .A1(g8068), .A2(g17262), .ZN(g19561) );
AND2_X4 U_g19562 ( .A1(g8076), .A2(g17265), .ZN(g19562) );
AND2_X4 U_g19564 ( .A1(g8123), .A2(g17272), .ZN(g19564) );
AND2_X4 U_g19565 ( .A1(g8126), .A2(g17275), .ZN(g19565) );
AND2_X4 U_g19566 ( .A1(g8129), .A2(g17278), .ZN(g19566) );
AND2_X4 U_g19567 ( .A1(g8138), .A2(g17282), .ZN(g19567) );
AND2_X4 U_g19568 ( .A1(g8141), .A2(g17285), .ZN(g19568) );
AND2_X4 U_g19569 ( .A1(g8144), .A2(g17288), .ZN(g19569) );
AND2_X4 U_g19570 ( .A1(g8150), .A2(g17291), .ZN(g19570) );
AND2_X4 U_g19571 ( .A1(g8153), .A2(g17294), .ZN(g19571) );
AND2_X4 U_g19572 ( .A1(g8161), .A2(g17297), .ZN(g19572) );
AND2_X4 U_g19574 ( .A1(g8191), .A2(g17304), .ZN(g19574) );
AND2_X4 U_g19575 ( .A1(g8194), .A2(g17307), .ZN(g19575) );
AND2_X4 U_g19576 ( .A1(g8197), .A2(g17310), .ZN(g19576) );
AND2_X4 U_g19584 ( .A1(g640), .A2(g18756), .ZN(g19584) );
AND2_X4 U_g19585 ( .A1(g692), .A2(g18757), .ZN(g19585) );
AND2_X4 U_g19586 ( .A1(g8209), .A2(g17315), .ZN(g19586) );
AND2_X4 U_g19587 ( .A1(g8212), .A2(g17318), .ZN(g19587) );
AND2_X4 U_g19588 ( .A1(g8215), .A2(g17321), .ZN(g19588) );
AND2_X4 U_g19589 ( .A1(g8224), .A2(g17324), .ZN(g19589) );
AND2_X4 U_g19590 ( .A1(g8227), .A2(g17327), .ZN(g19590) );
AND2_X4 U_g19591 ( .A1(g8230), .A2(g17330), .ZN(g19591) );
AND2_X4 U_g19592 ( .A1(g8236), .A2(g17333), .ZN(g19592) );
AND2_X4 U_g19593 ( .A1(g8239), .A2(g17336), .ZN(g19593) );
AND2_X4 U_g19594 ( .A1(g16935), .A2(g12555), .ZN(g19594) );
AND2_X4 U_g19597 ( .A1(g3922), .A2(g17342), .ZN(g19597) );
AND2_X4 U_g19598 ( .A1(g3925), .A2(g17345), .ZN(g19598) );
AND2_X4 U_g19599 ( .A1(g3928), .A2(g17348), .ZN(g19599) );
AND2_X4 U_g19600 ( .A1(g633), .A2(g18783), .ZN(g19600) );
AND2_X4 U_g19601 ( .A1(g640), .A2(g18784), .ZN(g19601) );
AND2_X4 U_g19602 ( .A1(g633), .A2(g18785), .ZN(g19602) );
AND2_X4 U_g19603 ( .A1(g692), .A2(g18786), .ZN(g19603) );
AND2_X4 U_g19604 ( .A1(g3948), .A2(g17354), .ZN(g19604) );
AND2_X4 U_g19605 ( .A1(g3951), .A2(g17357), .ZN(g19605) );
AND2_X4 U_g19606 ( .A1(g3954), .A2(g17360), .ZN(g19606) );
AND2_X4 U_g19614 ( .A1(g1326), .A2(g18787), .ZN(g19614) );
AND2_X4 U_g19615 ( .A1(g1378), .A2(g18788), .ZN(g19615) );
AND2_X4 U_g19616 ( .A1(g3966), .A2(g17363), .ZN(g19616) );
AND2_X4 U_g19617 ( .A1(g3969), .A2(g17366), .ZN(g19617) );
AND2_X4 U_g19618 ( .A1(g3972), .A2(g17369), .ZN(g19618) );
AND2_X4 U_g19619 ( .A1(g3981), .A2(g17372), .ZN(g19619) );
AND2_X4 U_g19620 ( .A1(g3984), .A2(g17375), .ZN(g19620) );
AND2_X4 U_g19621 ( .A1(g3987), .A2(g17378), .ZN(g19621) );
AND2_X4 U_g19623 ( .A1(g4000), .A2(g17384), .ZN(g19623) );
AND2_X4 U_g19624 ( .A1(g4003), .A2(g17387), .ZN(g19624) );
AND2_X4 U_g19625 ( .A1(g4006), .A2(g17390), .ZN(g19625) );
AND2_X4 U_g19626 ( .A1(g640), .A2(g18805), .ZN(g19626) );
AND2_X4 U_g19627 ( .A1(g633), .A2(g18806), .ZN(g19627) );
AND2_X4 U_g19628 ( .A1(g653), .A2(g18807), .ZN(g19628) );
AND2_X4 U_g19629 ( .A1(g692), .A2(g18808), .ZN(g19629) );
AND2_X4 U_g19630 ( .A1(g4029), .A2(g17399), .ZN(g19630) );
AND2_X4 U_g19631 ( .A1(g4032), .A2(g17402), .ZN(g19631) );
AND2_X4 U_g19632 ( .A1(g4035), .A2(g17405), .ZN(g19632) );
AND2_X4 U_g19633 ( .A1(g1319), .A2(g18809), .ZN(g19633) );
AND2_X4 U_g19634 ( .A1(g1326), .A2(g18810), .ZN(g19634) );
AND2_X4 U_g19635 ( .A1(g1319), .A2(g18811), .ZN(g19635) );
AND2_X4 U_g19636 ( .A1(g1378), .A2(g18812), .ZN(g19636) );
AND2_X4 U_g19637 ( .A1(g4055), .A2(g17410), .ZN(g19637) );
AND2_X4 U_g19638 ( .A1(g4058), .A2(g17413), .ZN(g19638) );
AND2_X4 U_g19639 ( .A1(g4061), .A2(g17416), .ZN(g19639) );
AND2_X4 U_g19647 ( .A1(g2020), .A2(g18813), .ZN(g19647) );
AND2_X4 U_g19648 ( .A1(g2072), .A2(g18814), .ZN(g19648) );
AND2_X4 U_g19649 ( .A1(g4073), .A2(g17419), .ZN(g19649) );
AND2_X4 U_g19650 ( .A1(g4076), .A2(g17422), .ZN(g19650) );
AND2_X4 U_g19651 ( .A1(g4079), .A2(g17425), .ZN(g19651) );
AND2_X4 U_g19653 ( .A1(g4095), .A2(g17430), .ZN(g19653) );
AND2_X4 U_g19654 ( .A1(g4098), .A2(g17433), .ZN(g19654) );
AND2_X4 U_g19655 ( .A1(g4101), .A2(g17436), .ZN(g19655) );
AND2_X4 U_g19656 ( .A1(g4104), .A2(g17439), .ZN(g19656) );
AND2_X4 U_g19660 ( .A1(g633), .A2(g18822), .ZN(g19660) );
AND2_X4 U_g19661 ( .A1(g653), .A2(g18823), .ZN(g19661) );
AND2_X4 U_g19662 ( .A1(g646), .A2(g18824), .ZN(g19662) );
AND2_X4 U_g19663 ( .A1(g4127), .A2(g17451), .ZN(g19663) );
AND2_X4 U_g19664 ( .A1(g4130), .A2(g17454), .ZN(g19664) );
AND2_X4 U_g19665 ( .A1(g4133), .A2(g17457), .ZN(g19665) );
AND2_X4 U_g19666 ( .A1(g1326), .A2(g18825), .ZN(g19666) );
AND2_X4 U_g19667 ( .A1(g1319), .A2(g18826), .ZN(g19667) );
AND2_X4 U_g19668 ( .A1(g1339), .A2(g18827), .ZN(g19668) );
AND2_X4 U_g19669 ( .A1(g1378), .A2(g18828), .ZN(g19669) );
AND2_X4 U_g19670 ( .A1(g4156), .A2(g17465), .ZN(g19670) );
AND2_X4 U_g19671 ( .A1(g4159), .A2(g17468), .ZN(g19671) );
AND2_X4 U_g19672 ( .A1(g4162), .A2(g17471), .ZN(g19672) );
AND2_X4 U_g19673 ( .A1(g2013), .A2(g18829), .ZN(g19673) );
AND2_X4 U_g19674 ( .A1(g2020), .A2(g18830), .ZN(g19674) );
AND2_X4 U_g19675 ( .A1(g2013), .A2(g18831), .ZN(g19675) );
AND2_X4 U_g19676 ( .A1(g2072), .A2(g18832), .ZN(g19676) );
AND2_X4 U_g19677 ( .A1(g4182), .A2(g17476), .ZN(g19677) );
AND2_X4 U_g19678 ( .A1(g4185), .A2(g17479), .ZN(g19678) );
AND2_X4 U_g19679 ( .A1(g4188), .A2(g17482), .ZN(g19679) );
AND2_X4 U_g19687 ( .A1(g2714), .A2(g18833), .ZN(g19687) );
AND2_X4 U_g19688 ( .A1(g2766), .A2(g18834), .ZN(g19688) );
AND2_X4 U_g19691 ( .A1(g16841), .A2(g10865), .ZN(g19691) );
AND2_X4 U_g19692 ( .A1(g4205), .A2(g17487), .ZN(g19692) );
AND2_X4 U_g19693 ( .A1(g4208), .A2(g17490), .ZN(g19693) );
AND2_X4 U_g19694 ( .A1(g4211), .A2(g17493), .ZN(g19694) );
AND2_X4 U_g19695 ( .A1(g4214), .A2(g17496), .ZN(g19695) );
AND2_X4 U_g19697 ( .A1(g653), .A2(g18838), .ZN(g19697) );
AND2_X4 U_g19698 ( .A1(g646), .A2(g18839), .ZN(g19698) );
AND2_X4 U_g19699 ( .A1(g660), .A2(g18840), .ZN(g19699) );
AND2_X4 U_g19700 ( .A1(g17815), .A2(g16024), .ZN(g19700) );
AND2_X4 U_g19701 ( .A1(g4234), .A2(g17511), .ZN(g19701) );
AND2_X4 U_g19702 ( .A1(g4237), .A2(g17514), .ZN(g19702) );
AND2_X4 U_g19703 ( .A1(g4240), .A2(g17517), .ZN(g19703) );
AND2_X4 U_g19704 ( .A1(g4243), .A2(g17520), .ZN(g19704) );
AND2_X4 U_g19708 ( .A1(g1319), .A2(g18841), .ZN(g19708) );
AND2_X4 U_g19709 ( .A1(g1339), .A2(g18842), .ZN(g19709) );
AND2_X4 U_g19710 ( .A1(g1332), .A2(g18843), .ZN(g19710) );
AND2_X4 U_g19711 ( .A1(g4266), .A2(g17531), .ZN(g19711) );
AND2_X4 U_g19712 ( .A1(g4269), .A2(g17534), .ZN(g19712) );
AND2_X4 U_g19713 ( .A1(g4272), .A2(g17537), .ZN(g19713) );
AND2_X4 U_g19714 ( .A1(g2020), .A2(g18844), .ZN(g19714) );
AND2_X4 U_g19715 ( .A1(g2013), .A2(g18845), .ZN(g19715) );
AND2_X4 U_g19716 ( .A1(g2033), .A2(g18846), .ZN(g19716) );
AND2_X4 U_g19717 ( .A1(g2072), .A2(g18847), .ZN(g19717) );
AND2_X4 U_g19718 ( .A1(g4295), .A2(g17545), .ZN(g19718) );
AND2_X4 U_g19719 ( .A1(g4298), .A2(g17548), .ZN(g19719) );
AND2_X4 U_g19720 ( .A1(g4301), .A2(g17551), .ZN(g19720) );
AND2_X4 U_g19721 ( .A1(g2707), .A2(g18848), .ZN(g19721) );
AND2_X4 U_g19722 ( .A1(g2714), .A2(g18849), .ZN(g19722) );
AND2_X4 U_g19723 ( .A1(g2707), .A2(g18850), .ZN(g19723) );
AND2_X4 U_g19724 ( .A1(g2766), .A2(g18851), .ZN(g19724) );
AND2_X4 U_g19726 ( .A1(g16847), .A2(g6131), .ZN(g19726) );
AND2_X4 U_g19727 ( .A1(g4329), .A2(g17557), .ZN(g19727) );
AND2_X4 U_g19728 ( .A1(g4332), .A2(g17560), .ZN(g19728) );
AND2_X4 U_g19729 ( .A1(g4335), .A2(g17563), .ZN(g19729) );
AND2_X4 U_g19730 ( .A1(g653), .A2(g17573), .ZN(g19730) );
AND2_X4 U_g19731 ( .A1(g646), .A2(g18853), .ZN(g19731) );
AND2_X4 U_g19732 ( .A1(g660), .A2(g18854), .ZN(g19732) );
AND2_X4 U_g19733 ( .A1(g672), .A2(g18855), .ZN(g19733) );
AND2_X4 U_g19734 ( .A1(g17815), .A2(g16034), .ZN(g19734) );
AND2_X4 U_g19735 ( .A1(g17903), .A2(g16035), .ZN(g19735) );
AND2_X4 U_g19736 ( .A1(g4360), .A2(g17579), .ZN(g19736) );
AND2_X4 U_g19737 ( .A1(g4363), .A2(g17582), .ZN(g19737) );
AND2_X4 U_g19738 ( .A1(g4366), .A2(g17585), .ZN(g19738) );
AND2_X4 U_g19739 ( .A1(g4369), .A2(g17588), .ZN(g19739) );
AND2_X4 U_g19741 ( .A1(g1339), .A2(g18856), .ZN(g19741) );
AND2_X4 U_g19742 ( .A1(g1332), .A2(g18857), .ZN(g19742) );
AND2_X4 U_g19743 ( .A1(g1346), .A2(g18858), .ZN(g19743) );
AND2_X4 U_g19744 ( .A1(g17927), .A2(g16040), .ZN(g19744) );
AND2_X4 U_g19745 ( .A1(g4389), .A2(g17601), .ZN(g19745) );
AND2_X4 U_g19746 ( .A1(g4392), .A2(g17604), .ZN(g19746) );
AND2_X4 U_g19747 ( .A1(g4395), .A2(g17607), .ZN(g19747) );
AND2_X4 U_g19748 ( .A1(g4398), .A2(g17610), .ZN(g19748) );
AND2_X4 U_g19752 ( .A1(g2013), .A2(g18859), .ZN(g19752) );
AND2_X4 U_g19753 ( .A1(g2033), .A2(g18860), .ZN(g19753) );
AND2_X4 U_g19754 ( .A1(g2026), .A2(g18861), .ZN(g19754) );
AND2_X4 U_g19755 ( .A1(g4421), .A2(g17621), .ZN(g19755) );
AND2_X4 U_g19756 ( .A1(g4424), .A2(g17624), .ZN(g19756) );
AND2_X4 U_g19757 ( .A1(g4427), .A2(g17627), .ZN(g19757) );
AND2_X4 U_g19758 ( .A1(g2714), .A2(g18862), .ZN(g19758) );
AND2_X4 U_g19759 ( .A1(g2707), .A2(g18863), .ZN(g19759) );
AND2_X4 U_g19760 ( .A1(g2727), .A2(g18864), .ZN(g19760) );
AND2_X4 U_g19761 ( .A1(g2766), .A2(g18865), .ZN(g19761) );
AND2_X4 U_g19764 ( .A1(g4453), .A2(g17637), .ZN(g19764) );
AND2_X4 U_g19765 ( .A1(g660), .A2(g18870), .ZN(g19765) );
AND2_X4 U_g19766 ( .A1(g672), .A2(g18871), .ZN(g19766) );
AND2_X4 U_g19767 ( .A1(g666), .A2(g18872), .ZN(g19767) );
AND2_X4 U_g19768 ( .A1(g17815), .A2(g16054), .ZN(g19768) );
AND2_X4 U_g19769 ( .A1(g17903), .A2(g16055), .ZN(g19769) );
AND2_X4 U_g19770 ( .A1(g4498), .A2(g17655), .ZN(g19770) );
AND2_X4 U_g19771 ( .A1(g4501), .A2(g17658), .ZN(g19771) );
AND2_X4 U_g19772 ( .A1(g4504), .A2(g17661), .ZN(g19772) );
AND2_X4 U_g19773 ( .A1(g1339), .A2(g17670), .ZN(g19773) );
AND2_X4 U_g19774 ( .A1(g1332), .A2(g18874), .ZN(g19774) );
AND2_X4 U_g19775 ( .A1(g1346), .A2(g18875), .ZN(g19775) );
AND2_X4 U_g19776 ( .A1(g1358), .A2(g18876), .ZN(g19776) );
AND2_X4 U_g19777 ( .A1(g17927), .A2(g16056), .ZN(g19777) );
AND2_X4 U_g19778 ( .A1(g18014), .A2(g16057), .ZN(g19778) );
AND2_X4 U_g19779 ( .A1(g4529), .A2(g17676), .ZN(g19779) );
AND2_X4 U_g19780 ( .A1(g4532), .A2(g17679), .ZN(g19780) );
AND2_X4 U_g19781 ( .A1(g4535), .A2(g17682), .ZN(g19781) );
AND2_X4 U_g19782 ( .A1(g4538), .A2(g17685), .ZN(g19782) );
AND2_X4 U_g19784 ( .A1(g2033), .A2(g18877), .ZN(g19784) );
AND2_X4 U_g19785 ( .A1(g2026), .A2(g18878), .ZN(g19785) );
AND2_X4 U_g19786 ( .A1(g2040), .A2(g18879), .ZN(g19786) );
AND2_X4 U_g19787 ( .A1(g18038), .A2(g16062), .ZN(g19787) );
AND2_X4 U_g19788 ( .A1(g4558), .A2(g17698), .ZN(g19788) );
AND2_X4 U_g19789 ( .A1(g4561), .A2(g17701), .ZN(g19789) );
AND2_X4 U_g19790 ( .A1(g4564), .A2(g17704), .ZN(g19790) );
AND2_X4 U_g19791 ( .A1(g4567), .A2(g17707), .ZN(g19791) );
AND2_X4 U_g19795 ( .A1(g2707), .A2(g18880), .ZN(g19795) );
AND2_X4 U_g19796 ( .A1(g2727), .A2(g18881), .ZN(g19796) );
AND2_X4 U_g19797 ( .A1(g2720), .A2(g18882), .ZN(g19797) );
AND3_X4 U_I26240 ( .A1(g18174), .A2(g18341), .A3(g17974), .ZN(I26240) );
AND3_X4 U_g19799 ( .A1(g17640), .A2(g18074), .A3(I26240), .ZN(g19799) );
AND2_X4 U_g19802 ( .A1(g672), .A2(g18891), .ZN(g19802) );
AND2_X4 U_g19803 ( .A1(g666), .A2(g18892), .ZN(g19803) );
AND2_X4 U_g19804 ( .A1(g679), .A2(g18893), .ZN(g19804) );
AND2_X4 U_g19805 ( .A1(g17903), .A2(g16088), .ZN(g19805) );
AND2_X4 U_g19806 ( .A1(g4629), .A2(g17738), .ZN(g19806) );
AND2_X4 U_g19807 ( .A1(g1346), .A2(g18896), .ZN(g19807) );
AND2_X4 U_g19808 ( .A1(g1358), .A2(g18897), .ZN(g19808) );
AND2_X4 U_g19809 ( .A1(g1352), .A2(g18898), .ZN(g19809) );
AND2_X4 U_g19810 ( .A1(g17927), .A2(g16090), .ZN(g19810) );
AND2_X4 U_g19811 ( .A1(g18014), .A2(g16091), .ZN(g19811) );
AND2_X4 U_g19812 ( .A1(g4674), .A2(g17755), .ZN(g19812) );
AND2_X4 U_g19813 ( .A1(g4677), .A2(g17758), .ZN(g19813) );
AND2_X4 U_g19814 ( .A1(g4680), .A2(g17761), .ZN(g19814) );
AND2_X4 U_g19815 ( .A1(g2033), .A2(g17770), .ZN(g19815) );
AND2_X4 U_g19816 ( .A1(g2026), .A2(g18900), .ZN(g19816) );
AND2_X4 U_g19817 ( .A1(g2040), .A2(g18901), .ZN(g19817) );
AND2_X4 U_g19818 ( .A1(g2052), .A2(g18902), .ZN(g19818) );
AND2_X4 U_g19819 ( .A1(g18038), .A2(g16092), .ZN(g19819) );
AND2_X4 U_g19820 ( .A1(g18131), .A2(g16093), .ZN(g19820) );
AND2_X4 U_g19821 ( .A1(g4705), .A2(g17776), .ZN(g19821) );
AND2_X4 U_g19822 ( .A1(g4708), .A2(g17779), .ZN(g19822) );
AND2_X4 U_g19823 ( .A1(g4711), .A2(g17782), .ZN(g19823) );
AND2_X4 U_g19824 ( .A1(g4714), .A2(g17785), .ZN(g19824) );
AND2_X4 U_g19826 ( .A1(g2727), .A2(g18903), .ZN(g19826) );
AND2_X4 U_g19827 ( .A1(g2720), .A2(g18904), .ZN(g19827) );
AND2_X4 U_g19828 ( .A1(g2734), .A2(g18905), .ZN(g19828) );
AND2_X4 U_g19829 ( .A1(g18155), .A2(g16098), .ZN(g19829) );
AND2_X4 U_g19836 ( .A1(g7143), .A2(g18908), .ZN(g19836) );
AND2_X4 U_g19837 ( .A1(g6901), .A2(g17799), .ZN(g19837) );
AND2_X4 U_g19839 ( .A1(g666), .A2(g18909), .ZN(g19839) );
AND2_X4 U_g19840 ( .A1(g679), .A2(g18910), .ZN(g19840) );
AND2_X4 U_g19841 ( .A1(g686), .A2(g18911), .ZN(g19841) );
AND3_X4 U_I26282 ( .A1(g18188), .A2(g18089), .A3(g17991), .ZN(I26282) );
AND3_X4 U_g19842 ( .A1(g14525), .A2(g13922), .A3(I26282), .ZN(g19842) );
AND3_X4 U_I26285 ( .A1(g18281), .A2(g18436), .A3(g18091), .ZN(I26285) );
AND3_X4 U_g19843 ( .A1(g17741), .A2(g18190), .A3(I26285), .ZN(g19843) );
AND2_X4 U_g19846 ( .A1(g1358), .A2(g18914), .ZN(g19846) );
AND2_X4 U_g19847 ( .A1(g1352), .A2(g18915), .ZN(g19847) );
AND2_X4 U_g19848 ( .A1(g1365), .A2(g18916), .ZN(g19848) );
AND2_X4 U_g19849 ( .A1(g18014), .A2(g16126), .ZN(g19849) );
AND2_X4 U_g19850 ( .A1(g4806), .A2(g17839), .ZN(g19850) );
AND2_X4 U_g19851 ( .A1(g2040), .A2(g18919), .ZN(g19851) );
AND2_X4 U_g19852 ( .A1(g2052), .A2(g18920), .ZN(g19852) );
AND2_X4 U_g19853 ( .A1(g2046), .A2(g18921), .ZN(g19853) );
AND2_X4 U_g19854 ( .A1(g18038), .A2(g16128), .ZN(g19854) );
AND2_X4 U_g19855 ( .A1(g18131), .A2(g16129), .ZN(g19855) );
AND2_X4 U_g19856 ( .A1(g4851), .A2(g17856), .ZN(g19856) );
AND2_X4 U_g19857 ( .A1(g4854), .A2(g17859), .ZN(g19857) );
AND2_X4 U_g19858 ( .A1(g4857), .A2(g17862), .ZN(g19858) );
AND2_X4 U_g19859 ( .A1(g2727), .A2(g17871), .ZN(g19859) );
AND2_X4 U_g19860 ( .A1(g2720), .A2(g18923), .ZN(g19860) );
AND2_X4 U_g19861 ( .A1(g2734), .A2(g18924), .ZN(g19861) );
AND2_X4 U_g19862 ( .A1(g2746), .A2(g18925), .ZN(g19862) );
AND2_X4 U_g19863 ( .A1(g18155), .A2(g16130), .ZN(g19863) );
AND2_X4 U_g19864 ( .A1(g18247), .A2(g16131), .ZN(g19864) );
AND3_X4 U_g19868 ( .A1(g16498), .A2(g16867), .A3(g19001), .ZN(g19868) );
AND2_X4 U_g19869 ( .A1(g679), .A2(g18926), .ZN(g19869) );
AND2_X4 U_g19870 ( .A1(g686), .A2(g18927), .ZN(g19870) );
AND3_X4 U_I26311 ( .A1(g18353), .A2(g13958), .A3(g14011), .ZN(I26311) );
AND3_X4 U_g19871 ( .A1(g14086), .A2(g18275), .A3(I26311), .ZN(g19871) );
AND2_X4 U_g19872 ( .A1(g1352), .A2(g18928), .ZN(g19872) );
AND2_X4 U_g19873 ( .A1(g1365), .A2(g18929), .ZN(g19873) );
AND2_X4 U_g19874 ( .A1(g1372), .A2(g18930), .ZN(g19874) );
AND3_X4 U_I26317 ( .A1(g18295), .A2(g18205), .A3(g18108), .ZN(I26317) );
AND3_X4 U_g19875 ( .A1(g14580), .A2(g13978), .A3(I26317), .ZN(g19875) );
AND3_X4 U_I26320 ( .A1(g18374), .A2(g18509), .A3(g18207), .ZN(I26320) );
AND3_X4 U_g19876 ( .A1(g17842), .A2(g18297), .A3(I26320), .ZN(g19876) );
AND2_X4 U_g19879 ( .A1(g2052), .A2(g18933), .ZN(g19879) );
AND2_X4 U_g19880 ( .A1(g2046), .A2(g18934), .ZN(g19880) );
AND2_X4 U_g19881 ( .A1(g2059), .A2(g18935), .ZN(g19881) );
AND2_X4 U_g19882 ( .A1(g18131), .A2(g16177), .ZN(g19882) );
AND2_X4 U_g19883 ( .A1(g4982), .A2(g17951), .ZN(g19883) );
AND2_X4 U_g19884 ( .A1(g2734), .A2(g18938), .ZN(g19884) );
AND2_X4 U_g19885 ( .A1(g2746), .A2(g18939), .ZN(g19885) );
AND2_X4 U_g19886 ( .A1(g2740), .A2(g18940), .ZN(g19886) );
AND2_X4 U_g19887 ( .A1(g18155), .A2(g16179), .ZN(g19887) );
AND2_X4 U_g19888 ( .A1(g18247), .A2(g16180), .ZN(g19888) );
AND2_X4 U_g19889 ( .A1(g2912), .A2(g18943), .ZN(g19889) );
AND2_X4 U_g19895 ( .A1(g686), .A2(g18945), .ZN(g19895) );
AND3_X4 U_g19899 ( .A1(g16520), .A2(g16895), .A3(g16507), .ZN(g19899) );
AND2_X4 U_g19900 ( .A1(g1365), .A2(g18946), .ZN(g19900) );
AND2_X4 U_g19901 ( .A1(g1372), .A2(g18947), .ZN(g19901) );
AND3_X4 U_I26348 ( .A1(g18448), .A2(g14028), .A3(g14102), .ZN(I26348) );
AND3_X4 U_g19902 ( .A1(g14201), .A2(g18368), .A3(I26348), .ZN(g19902) );
AND2_X4 U_g19903 ( .A1(g2046), .A2(g18948), .ZN(g19903) );
AND2_X4 U_g19904 ( .A1(g2059), .A2(g18949), .ZN(g19904) );
AND2_X4 U_g19905 ( .A1(g2066), .A2(g18950), .ZN(g19905) );
AND3_X4 U_I26354 ( .A1(g18388), .A2(g18312), .A3(g18224), .ZN(I26354) );
AND3_X4 U_g19906 ( .A1(g14614), .A2(g14048), .A3(I26354), .ZN(g19906) );
AND3_X4 U_I26357 ( .A1(g18469), .A2(g18573), .A3(g18314), .ZN(I26357) );
AND3_X4 U_g19907 ( .A1(g17954), .A2(g18390), .A3(I26357), .ZN(g19907) );
AND2_X4 U_g19910 ( .A1(g2746), .A2(g18953), .ZN(g19910) );
AND2_X4 U_g19911 ( .A1(g2740), .A2(g18954), .ZN(g19911) );
AND2_X4 U_g19912 ( .A1(g2753), .A2(g18955), .ZN(g19912) );
AND2_X4 U_g19913 ( .A1(g18247), .A2(g16236), .ZN(g19913) );
AND2_X4 U_g19914 ( .A1(g3018), .A2(g18958), .ZN(g19914) );
AND2_X4 U_g19920 ( .A1(g1372), .A2(g18961), .ZN(g19920) );
AND3_X4 U_g19924 ( .A1(g16551), .A2(g16924), .A3(g16529), .ZN(g19924) );
AND2_X4 U_g19925 ( .A1(g2059), .A2(g18962), .ZN(g19925) );
AND2_X4 U_g19926 ( .A1(g2066), .A2(g18963), .ZN(g19926) );
AND3_X4 U_I26377 ( .A1(g18521), .A2(g14119), .A3(g14217), .ZN(I26377) );
AND3_X4 U_g19927 ( .A1(g14316), .A2(g18463), .A3(I26377), .ZN(g19927) );
AND2_X4 U_g19928 ( .A1(g2740), .A2(g18964), .ZN(g19928) );
AND2_X4 U_g19929 ( .A1(g2753), .A2(g18965), .ZN(g19929) );
AND2_X4 U_g19930 ( .A1(g2760), .A2(g18966), .ZN(g19930) );
AND3_X4 U_I26383 ( .A1(g18483), .A2(g18405), .A3(g18331), .ZN(I26383) );
AND3_X4 U_g19931 ( .A1(g14637), .A2(g14139), .A3(I26383), .ZN(g19931) );
AND2_X4 U_g19932 ( .A1(g2917), .A2(g18166), .ZN(g19932) );
AND2_X4 U_g19935 ( .A1(g2066), .A2(g18972), .ZN(g19935) );
AND3_X4 U_g19939 ( .A1(g16583), .A2(g16954), .A3(g16560), .ZN(g19939) );
AND2_X4 U_g19940 ( .A1(g2753), .A2(g18973), .ZN(g19940) );
AND2_X4 U_g19941 ( .A1(g2760), .A2(g18974), .ZN(g19941) );
AND3_X4 U_I26396 ( .A1(g18585), .A2(g14234), .A3(g14332), .ZN(I26396) );
AND3_X4 U_g19942 ( .A1(g14438), .A2(g18536), .A3(I26396), .ZN(g19942) );
AND2_X4 U_g19943 ( .A1(g7562), .A2(g18976), .ZN(g19943) );
AND2_X4 U_g19944 ( .A1(g3028), .A2(g18258), .ZN(g19944) );
AND2_X4 U_g19949 ( .A1(g5293), .A2(g18278), .ZN(g19949) );
AND2_X4 U_g19952 ( .A1(g2760), .A2(g18987), .ZN(g19952) );
AND2_X4 U_g19953 ( .A1(g7566), .A2(g18334), .ZN(g19953) );
AND3_X4 U_I26416 ( .A1(g18553), .A2(g18491), .A3(g18431), .ZN(I26416) );
AND3_X4 U_g19970 ( .A1(g18354), .A2(g18276), .A3(I26416), .ZN(g19970) );
AND2_X4 U_g19971 ( .A1(g5327), .A2(g18355), .ZN(g19971) );
AND2_X4 U_g19976 ( .A1(g5330), .A2(g18371), .ZN(g19976) );
AND3_X4 U_I26432 ( .A1(g18277), .A2(g18189), .A3(g18090), .ZN(I26432) );
AND3_X4 U_g19982 ( .A1(g17992), .A2(g17913), .A3(I26432), .ZN(g19982) );
AND2_X4 U_g19983 ( .A1(g5352), .A2(g18432), .ZN(g19983) );
AND3_X4 U_I26440 ( .A1(g18603), .A2(g18555), .A3(g18504), .ZN(I26440) );
AND3_X4 U_g20000 ( .A1(g18449), .A2(g18369), .A3(I26440), .ZN(g20000) );
AND2_X4 U_g20001 ( .A1(g5355), .A2(g18450), .ZN(g20001) );
AND2_X4 U_g20006 ( .A1(g5358), .A2(g18466), .ZN(g20006) );
AND2_X4 U_g20011 ( .A1(g18063), .A2(g3113), .ZN(g20011) );
AND2_X4 U_g20012 ( .A1(g16804), .A2(g3135), .ZN(g20012) );
AND2_X4 U_g20013 ( .A1(g17720), .A2(g12848), .ZN(g20013) );
AND2_X4 U_g20014 ( .A1(g7615), .A2(g16749), .ZN(g20014) );
AND3_X4 U_I26464 ( .A1(g18370), .A2(g18296), .A3(g18206), .ZN(I26464) );
AND3_X4 U_g20020 ( .A1(g18109), .A2(g18024), .A3(I26464), .ZN(g20020) );
AND2_X4 U_g20021 ( .A1(g5369), .A2(g18505), .ZN(g20021) );
AND3_X4 U_I26472 ( .A1(g18635), .A2(g18605), .A3(g18568), .ZN(I26472) );
AND3_X4 U_g20038 ( .A1(g18522), .A2(g18464), .A3(I26472), .ZN(g20038) );
AND2_X4 U_g20039 ( .A1(g5372), .A2(g18523), .ZN(g20039) );
AND2_X4 U_g20044 ( .A1(g5375), .A2(g18539), .ZN(g20044) );
AND2_X4 U_g20048 ( .A1(g16749), .A2(g3127), .ZN(g20048) );
AND2_X4 U_g20049 ( .A1(g17878), .A2(g3155), .ZN(g20049) );
AND2_X4 U_g20050 ( .A1(g18070), .A2(g3161), .ZN(g20050) );
AND2_X4 U_g20051 ( .A1(g18063), .A2(g3114), .ZN(g20051) );
AND2_X4 U_g20052 ( .A1(g16804), .A2(g3134), .ZN(g20052) );
AND2_X4 U_g20053 ( .A1(g17720), .A2(g12875), .ZN(g20053) );
AND3_X4 U_I26500 ( .A1(g18465), .A2(g18389), .A3(g18313), .ZN(I26500) );
AND3_X4 U_g20062 ( .A1(g18225), .A2(g18141), .A3(I26500), .ZN(g20062) );
AND2_X4 U_g20063 ( .A1(g5382), .A2(g18569), .ZN(g20063) );
AND3_X4 U_I26508 ( .A1(g18644), .A2(g18637), .A3(g18618), .ZN(I26508) );
AND3_X4 U_g20080 ( .A1(g18586), .A2(g18537), .A3(I26508), .ZN(g20080) );
AND2_X4 U_g20081 ( .A1(g5385), .A2(g18587), .ZN(g20081) );
AND2_X4 U_g20084 ( .A1(g17969), .A2(g3158), .ZN(g20084) );
AND2_X4 U_g20085 ( .A1(g18170), .A2(g3164), .ZN(g20085) );
AND2_X4 U_g20086 ( .A1(g18337), .A2(g3170), .ZN(g20086) );
AND2_X4 U_g20087 ( .A1(g16749), .A2(g7574), .ZN(g20087) );
AND2_X4 U_g20088 ( .A1(g16836), .A2(g3147), .ZN(g20088) );
AND2_X4 U_g20089 ( .A1(g17969), .A2(g9160), .ZN(g20089) );
AND2_X4 U_g20090 ( .A1(g18063), .A2(g3120), .ZN(g20090) );
AND2_X4 U_g20091 ( .A1(g16804), .A2(g3136), .ZN(g20091) );
AND2_X4 U_g20092 ( .A1(g16749), .A2(g7603), .ZN(g20092) );
AND3_X4 U_I26525 ( .A1(g18656), .A2(g18670), .A3(g18692), .ZN(I26525) );
AND4_X4 U_g20093 ( .A1(g13657), .A2(g13677), .A3(g13750), .A4(I26525), .ZN(g20093) );
AND3_X4 U_I26528 ( .A1(g18656), .A2(g14837), .A3(g13657), .ZN(I26528) );
AND3_X4 U_g20094 ( .A1(g13677), .A2(g13706), .A3(I26528), .ZN(g20094) );
AND3_X4 U_I26541 ( .A1(g18538), .A2(g18484), .A3(g18406), .ZN(I26541) );
AND3_X4 U_g20103 ( .A1(g18332), .A2(g18257), .A3(I26541), .ZN(g20103) );
AND2_X4 U_g20104 ( .A1(g5391), .A2(g18619), .ZN(g20104) );
AND2_X4 U_g20106 ( .A1(g18261), .A2(g3167), .ZN(g20106) );
AND2_X4 U_g20107 ( .A1(g18415), .A2(g3173), .ZN(g20107) );
AND2_X4 U_g20108 ( .A1(g18543), .A2(g3179), .ZN(g20108) );
AND2_X4 U_g20109 ( .A1(g17878), .A2(g9504), .ZN(g20109) );
AND2_X4 U_g20110 ( .A1(g18070), .A2(g9286), .ZN(g20110) );
AND2_X4 U_g20111 ( .A1(g18261), .A2(g9884), .ZN(g20111) );
AND2_X4 U_g20112 ( .A1(g16749), .A2(g3132), .ZN(g20112) );
AND2_X4 U_g20113 ( .A1(g16836), .A2(g3142), .ZN(g20113) );
AND2_X4 U_g20114 ( .A1(g17969), .A2(g9755), .ZN(g20114) );
AND2_X4 U_g20115 ( .A1(g16804), .A2(g3139), .ZN(g20115) );
AND3_X4 U_I26558 ( .A1(g14776), .A2(g18670), .A3(g18720), .ZN(I26558) );
AND4_X4 U_g20116 ( .A1(g16142), .A2(g13677), .A3(g13706), .A4(I26558), .ZN(g20116) );
AND3_X4 U_I26561 ( .A1(g14776), .A2(g18720), .A3(g13657), .ZN(I26561) );
AND3_X4 U_g20117 ( .A1(g16189), .A2(g13706), .A3(I26561), .ZN(g20117) );
AND3_X4 U_I26564 ( .A1(g18679), .A2(g18699), .A3(g18728), .ZN(I26564) );
AND4_X4 U_g20118 ( .A1(g13687), .A2(g13714), .A3(g13791), .A4(I26564), .ZN(g20118) );
AND3_X4 U_I26567 ( .A1(g18679), .A2(g14910), .A3(g13687), .ZN(I26567) );
AND3_X4 U_g20119 ( .A1(g13714), .A2(g13756), .A3(I26567), .ZN(g20119) );
AND2_X4 U_g20131 ( .A1(g18486), .A2(g3176), .ZN(g20131) );
AND2_X4 U_g20132 ( .A1(g18593), .A2(g3182), .ZN(g20132) );
AND2_X4 U_g20133 ( .A1(g18170), .A2(g9505), .ZN(g20133) );
AND2_X4 U_g20134 ( .A1(g18337), .A2(g9506), .ZN(g20134) );
AND2_X4 U_g20135 ( .A1(g18486), .A2(g9885), .ZN(g20135) );
AND2_X4 U_g20136 ( .A1(g17878), .A2(g9423), .ZN(g20136) );
AND2_X4 U_g20137 ( .A1(g18070), .A2(g9226), .ZN(g20137) );
AND2_X4 U_g20138 ( .A1(g18261), .A2(g9756), .ZN(g20138) );
AND2_X4 U_g20139 ( .A1(g16836), .A2(g3151), .ZN(g20139) );
AND3_X4 U_g20144 ( .A1(g16679), .A2(g16884), .A3(g16665), .ZN(g20144) );
AND4_X4 U_g20145 ( .A1(g14776), .A2(g18670), .A3(g16142), .A4(g16189), .ZN(g20145) );
AND3_X4 U_I26590 ( .A1(g14811), .A2(g18699), .A3(g18758), .ZN(I26590) );
AND4_X4 U_g20146 ( .A1(g16201), .A2(g13714), .A3(g13756), .A4(I26590), .ZN(g20146) );
AND3_X4 U_I26593 ( .A1(g14811), .A2(g18758), .A3(g13687), .ZN(I26593) );
AND3_X4 U_g20147 ( .A1(g16254), .A2(g13756), .A3(I26593), .ZN(g20147) );
AND3_X4 U_I26596 ( .A1(g18708), .A2(g18735), .A3(g18765), .ZN(I26596) );
AND4_X4 U_g20148 ( .A1(g13724), .A2(g13764), .A3(g13819), .A4(I26596), .ZN(g20148) );
AND3_X4 U_I26599 ( .A1(g18708), .A2(g14991), .A3(g13724), .ZN(I26599) );
AND3_X4 U_g20149 ( .A1(g13764), .A2(g13797), .A3(I26599), .ZN(g20149) );
AND2_X4 U_g20156 ( .A1(g16809), .A2(g3185), .ZN(g20156) );
AND2_X4 U_g20157 ( .A1(g18415), .A2(g9287), .ZN(g20157) );
AND2_X4 U_g20158 ( .A1(g18543), .A2(g9886), .ZN(g20158) );
AND2_X4 U_g20159 ( .A1(g16809), .A2(g9288), .ZN(g20159) );
AND2_X4 U_g20160 ( .A1(g18170), .A2(g9424), .ZN(g20160) );
AND2_X4 U_g20161 ( .A1(g18337), .A2(g9426), .ZN(g20161) );
AND2_X4 U_g20162 ( .A1(g18486), .A2(g9757), .ZN(g20162) );
AND3_X4 U_I26615 ( .A1(g14797), .A2(g18692), .A3(g13657), .ZN(I26615) );
AND3_X4 U_g20177 ( .A1(g13677), .A2(g13750), .A3(I26615), .ZN(g20177) );
AND3_X4 U_g20182 ( .A1(g16705), .A2(g16913), .A3(g16686), .ZN(g20182) );
AND4_X4 U_g20183 ( .A1(g14811), .A2(g18699), .A3(g16201), .A4(g16254), .ZN(g20183) );
AND3_X4 U_I26621 ( .A1(g14863), .A2(g18735), .A3(g18789), .ZN(I26621) );
AND4_X4 U_g20184 ( .A1(g16266), .A2(g13764), .A3(g13797), .A4(I26621), .ZN(g20184) );
AND3_X4 U_I26624 ( .A1(g14863), .A2(g18789), .A3(g13724), .ZN(I26624) );
AND3_X4 U_g20185 ( .A1(g16313), .A2(g13797), .A3(I26624), .ZN(g20185) );
AND3_X4 U_I26627 ( .A1(g18744), .A2(g18772), .A3(g18796), .ZN(I26627) );
AND4_X4 U_g20186 ( .A1(g13774), .A2(g13805), .A3(g13840), .A4(I26627), .ZN(g20186) );
AND3_X4 U_I26630 ( .A1(g18744), .A2(g15080), .A3(g13774), .ZN(I26630) );
AND3_X4 U_g20187 ( .A1(g13805), .A2(g13825), .A3(I26630), .ZN(g20187) );
AND2_X4 U_g20188 ( .A1(g18593), .A2(g9425), .ZN(g20188) );
AND2_X4 U_g20189 ( .A1(g16825), .A2(g9289), .ZN(g20189) );
AND2_X4 U_g20190 ( .A1(g18415), .A2(g9227), .ZN(g20190) );
AND2_X4 U_g20191 ( .A1(g18543), .A2(g9758), .ZN(g20191) );
AND2_X4 U_g20192 ( .A1(g16809), .A2(g9228), .ZN(g20192) );
AND3_X4 U_I26639 ( .A1(g18656), .A2(g18670), .A3(g16142), .ZN(I26639) );
AND3_X4 U_g20197 ( .A1(g13677), .A2(g13706), .A3(I26639), .ZN(g20197) );
AND3_X4 U_I26645 ( .A1(g14849), .A2(g18728), .A3(g13687), .ZN(I26645) );
AND3_X4 U_g20211 ( .A1(g13714), .A2(g13791), .A3(I26645), .ZN(g20211) );
AND3_X4 U_g20216 ( .A1(g16736), .A2(g16943), .A3(g16712), .ZN(g20216) );
AND4_X4 U_g20217 ( .A1(g14863), .A2(g18735), .A3(g16266), .A4(g16313), .ZN(g20217) );
AND3_X4 U_I26651 ( .A1(g14936), .A2(g18772), .A3(g18815), .ZN(I26651) );
AND4_X4 U_g20218 ( .A1(g16325), .A2(g13805), .A3(g13825), .A4(I26651), .ZN(g20218) );
AND3_X4 U_I26654 ( .A1(g14936), .A2(g18815), .A3(g13774), .ZN(I26654) );
AND3_X4 U_g20219 ( .A1(g16371), .A2(g13825), .A3(I26654), .ZN(g20219) );
AND2_X4 U_g20220 ( .A1(g18593), .A2(g9355), .ZN(g20220) );
AND2_X4 U_g20221 ( .A1(g16825), .A2(g10099), .ZN(g20221) );
AND4_X4 U_g20222 ( .A1(g18656), .A2(g18720), .A3(g13657), .A4(g16293), .ZN(g20222) );
AND3_X4 U_I26661 ( .A1(g18679), .A2(g18699), .A3(g16201), .ZN(I26661) );
AND3_X4 U_g20227 ( .A1(g13714), .A2(g13756), .A3(I26661), .ZN(g20227) );
AND3_X4 U_I26667 ( .A1(g14922), .A2(g18765), .A3(g13724), .ZN(I26667) );
AND3_X4 U_g20241 ( .A1(g13764), .A2(g13819), .A3(I26667), .ZN(g20241) );
AND3_X4 U_g20246 ( .A1(g16778), .A2(g16974), .A3(g16743), .ZN(g20246) );
AND4_X4 U_g20247 ( .A1(g14936), .A2(g18772), .A3(g16325), .A4(g16371), .ZN(g20247) );
AND3_X4 U_g20248 ( .A1(g18656), .A2(g14837), .A3(g16293), .ZN(g20248) );
AND4_X4 U_g20249 ( .A1(g18679), .A2(g18758), .A3(g13687), .A4(g16351), .ZN(g20249) );
AND3_X4 U_I26676 ( .A1(g18708), .A2(g18735), .A3(g16266), .ZN(I26676) );
AND3_X4 U_g20254 ( .A1(g13764), .A2(g13797), .A3(I26676), .ZN(g20254) );
AND3_X4 U_I26682 ( .A1(g15003), .A2(g18796), .A3(g13774), .ZN(I26682) );
AND3_X4 U_g20268 ( .A1(g13805), .A2(g13840), .A3(I26682), .ZN(g20268) );
AND4_X4 U_g20270 ( .A1(g14797), .A2(g18692), .A3(g13657), .A4(g16243), .ZN(g20270) );
AND3_X4 U_g20271 ( .A1(g18679), .A2(g14910), .A3(g16351), .ZN(g20271) );
AND4_X4 U_g20272 ( .A1(g18708), .A2(g18789), .A3(g13724), .A4(g16395), .ZN(g20272) );
AND3_X4 U_I26690 ( .A1(g18744), .A2(g18772), .A3(g16325), .ZN(I26690) );
AND3_X4 U_g20277 ( .A1(g13805), .A2(g13825), .A3(I26690), .ZN(g20277) );
AND3_X4 U_I26695 ( .A1(g18670), .A2(g18692), .A3(g16142), .ZN(I26695) );
AND3_X4 U_g20280 ( .A1(g13677), .A2(g16243), .A3(I26695), .ZN(g20280) );
AND4_X4 U_g20282 ( .A1(g14849), .A2(g18728), .A3(g13687), .A4(g16302), .ZN(g20282) );
AND3_X4 U_g20283 ( .A1(g18708), .A2(g14991), .A3(g16395), .ZN(g20283) );
AND4_X4 U_g20284 ( .A1(g18744), .A2(g18815), .A3(g13774), .A4(g16433), .ZN(g20284) );
AND2_X4 U_g20285 ( .A1(g16846), .A2(g8103), .ZN(g20285) );
AND3_X4 U_I26708 ( .A1(g18699), .A2(g18728), .A3(g16201), .ZN(I26708) );
AND3_X4 U_g20291 ( .A1(g13714), .A2(g16302), .A3(I26708), .ZN(g20291) );
AND4_X4 U_g20293 ( .A1(g14922), .A2(g18765), .A3(g13724), .A4(g16360), .ZN(g20293) );
AND3_X4 U_g20294 ( .A1(g18744), .A2(g15080), .A3(g16433), .ZN(g20294) );
AND3_X4 U_I26726 ( .A1(g18735), .A2(g18765), .A3(g16266), .ZN(I26726) );
AND3_X4 U_g20307 ( .A1(g13764), .A2(g16360), .A3(I26726), .ZN(g20307) );
AND4_X4 U_g20309 ( .A1(g15003), .A2(g18796), .A3(g13774), .A4(g16404), .ZN(g20309) );
AND3_X4 U_I26745 ( .A1(g18772), .A2(g18796), .A3(g16325), .ZN(I26745) );
AND3_X4 U_g20326 ( .A1(g13805), .A2(g16404), .A3(I26745), .ZN(g20326) );
AND2_X4 U_g20460 ( .A1(g17351), .A2(g13644), .ZN(g20460) );
AND2_X4 U_g20472 ( .A1(g17314), .A2(g13669), .ZN(g20472) );
AND2_X4 U_g20480 ( .A1(g17313), .A2(g11827), .ZN(g20480) );
AND2_X4 U_g20486 ( .A1(g17281), .A2(g11859), .ZN(g20486) );
AND2_X4 U_g20492 ( .A1(g17258), .A2(g11894), .ZN(g20492) );
AND2_X4 U_g20499 ( .A1(g17648), .A2(g11933), .ZN(g20499) );
AND2_X4 U_g20502 ( .A1(g17566), .A2(g11973), .ZN(g20502) );
AND2_X4 U_g20503 ( .A1(g17507), .A2(g13817), .ZN(g20503) );
AND2_X4 U_g20506 ( .A1(g17499), .A2(g12025), .ZN(g20506) );
AND2_X4 U_g20512 ( .A1(g17445), .A2(g13836), .ZN(g20512) );
AND2_X4 U_g20525 ( .A1(g17394), .A2(g13849), .ZN(g20525) );
AND4_X4 U_g20538 ( .A1(g18656), .A2(g14837), .A3(g13657), .A4(g16189), .ZN(g20538) );
AND2_X4 U_g20640 ( .A1(g4809), .A2(g19064), .ZN(g20640) );
AND2_X4 U_g20647 ( .A1(g5888), .A2(g19075), .ZN(g20647) );
AND2_X4 U_g20665 ( .A1(g4985), .A2(g19081), .ZN(g20665) );
AND2_X4 U_g20809 ( .A1(g5712), .A2(g19113), .ZN(g20809) );
AND2_X4 U_g20826 ( .A1(g5770), .A2(g19118), .ZN(g20826) );
AND2_X4 U_g20836 ( .A1(g5829), .A2(g19125), .ZN(g20836) );
AND2_X4 U_g20840 ( .A1(g5885), .A2(g19132), .ZN(g20840) );
AND3_X4 U_g21049 ( .A1(g20016), .A2(g14079), .A3(g14165), .ZN(g21049) );
AND2_X4 U_g21067 ( .A1(g20193), .A2(g12030), .ZN(g21067) );
AND3_X4 U_g21068 ( .A1(g20058), .A2(g14194), .A3(g14280), .ZN(g21068) );
AND2_X4 U_g21077 ( .A1(g20223), .A2(g12094), .ZN(g21077) );
AND3_X4 U_g21078 ( .A1(g20099), .A2(g14309), .A3(g14402), .ZN(g21078) );
AND3_X4 U_g21085 ( .A1(g19484), .A2(g14158), .A3(g19001), .ZN(g21085) );
AND2_X4 U_g21086 ( .A1(g20193), .A2(g12142), .ZN(g21086) );
AND2_X4 U_g21091 ( .A1(g20250), .A2(g12166), .ZN(g21091) );
AND3_X4 U_g21092 ( .A1(g20124), .A2(g14431), .A3(g14514), .ZN(g21092) );
AND3_X4 U_g21097 ( .A1(g19505), .A2(g14273), .A3(g16507), .ZN(g21097) );
AND2_X4 U_g21098 ( .A1(g20223), .A2(g12204), .ZN(g21098) );
AND2_X4 U_g21103 ( .A1(g20273), .A2(g12228), .ZN(g21103) );
AND3_X4 U_g21107 ( .A1(g19444), .A2(g17893), .A3(g14079), .ZN(g21107) );
AND3_X4 U_g21111 ( .A1(g19524), .A2(g14395), .A3(g16529), .ZN(g21111) );
AND2_X4 U_g21112 ( .A1(g20250), .A2(g12259), .ZN(g21112) );
AND2_X4 U_g21121 ( .A1(g20054), .A2(g14244), .ZN(g21121) );
AND2_X4 U_g21122 ( .A1(g20140), .A2(g12279), .ZN(g21122) );
AND2_X4 U_g21123 ( .A1(g19970), .A2(g19982), .ZN(g21123) );
AND3_X4 U_g21124 ( .A1(g19471), .A2(g18004), .A3(g14194), .ZN(g21124) );
AND3_X4 U_g21128 ( .A1(g19534), .A2(g14507), .A3(g16560), .ZN(g21128) );
AND2_X4 U_g21129 ( .A1(g20273), .A2(g12302), .ZN(g21129) );
AND3_X4 U_I27695 ( .A1(g19318), .A2(g19300), .A3(g19286), .ZN(I27695) );
AND3_X4 U_g21136 ( .A1(g19271), .A2(g19261), .A3(I27695), .ZN(g21136) );
AND2_X4 U_g21137 ( .A1(g5750), .A2(g19272), .ZN(g21137) );
AND2_X4 U_g21138 ( .A1(g19484), .A2(g14347), .ZN(g21138) );
AND2_X4 U_g21140 ( .A1(g20095), .A2(g14366), .ZN(g21140) );
AND2_X4 U_g21141 ( .A1(g20178), .A2(g12315), .ZN(g21141) );
AND2_X4 U_g21142 ( .A1(g20000), .A2(g20020), .ZN(g21142) );
AND3_X4 U_g21143 ( .A1(g19494), .A2(g18121), .A3(g14309), .ZN(g21143) );
AND3_X4 U_I27711 ( .A1(g19262), .A2(g19414), .A3(g19386), .ZN(I27711) );
AND3_X4 U_g21152 ( .A1(g19357), .A2(g19334), .A3(I27711), .ZN(g21152) );
AND3_X4 U_g21153 ( .A1(g20054), .A2(g16543), .A3(g16501), .ZN(g21153) );
AND2_X4 U_g21154 ( .A1(g20193), .A2(g12333), .ZN(g21154) );
AND2_X4 U_g21155 ( .A1(g20140), .A2(g12336), .ZN(g21155) );
AND3_X4 U_I27717 ( .A1(g19345), .A2(g19321), .A3(g19304), .ZN(I27717) );
AND3_X4 U_g21156 ( .A1(g19290), .A2(g19276), .A3(I27717), .ZN(g21156) );
AND2_X4 U_g21157 ( .A1(g5809), .A2(g19291), .ZN(g21157) );
AND2_X4 U_g21158 ( .A1(g19505), .A2(g14459), .ZN(g21158) );
AND2_X4 U_g21160 ( .A1(g20120), .A2(g14478), .ZN(g21160) );
AND2_X4 U_g21161 ( .A1(g20212), .A2(g12343), .ZN(g21161) );
AND2_X4 U_g21162 ( .A1(g20038), .A2(g20062), .ZN(g21162) );
AND3_X4 U_g21163 ( .A1(g19515), .A2(g18237), .A3(g14431), .ZN(g21163) );
AND3_X4 U_I27733 ( .A1(g19277), .A2(g19451), .A3(g19416), .ZN(I27733) );
AND3_X4 U_g21172 ( .A1(g19389), .A2(g19368), .A3(I27733), .ZN(g21172) );
AND3_X4 U_g21173 ( .A1(g20095), .A2(g16575), .A3(g16523), .ZN(g21173) );
AND2_X4 U_g21174 ( .A1(g20223), .A2(g12363), .ZN(g21174) );
AND2_X4 U_g21175 ( .A1(g20178), .A2(g12366), .ZN(g21175) );
AND3_X4 U_I27739 ( .A1(g19379), .A2(g19348), .A3(g19325), .ZN(I27739) );
AND3_X4 U_g21176 ( .A1(g19308), .A2(g19295), .A3(I27739), .ZN(g21176) );
AND2_X4 U_g21177 ( .A1(g5865), .A2(g19309), .ZN(g21177) );
AND2_X4 U_g21178 ( .A1(g19524), .A2(g14546), .ZN(g21178) );
AND2_X4 U_g21180 ( .A1(g20150), .A2(g14565), .ZN(g21180) );
AND2_X4 U_g21181 ( .A1(g20242), .A2(g12373), .ZN(g21181) );
AND2_X4 U_g21182 ( .A1(g20080), .A2(g20103), .ZN(g21182) );
AND2_X4 U_g21188 ( .A1(g20140), .A2(g12379), .ZN(g21188) );
AND3_X4 U_I27755 ( .A1(g19296), .A2(g19478), .A3(g19453), .ZN(I27755) );
AND3_X4 U_g21192 ( .A1(g19419), .A2(g19400), .A3(I27755), .ZN(g21192) );
AND3_X4 U_g21193 ( .A1(g20120), .A2(g16599), .A3(g16554), .ZN(g21193) );
AND2_X4 U_g21194 ( .A1(g20250), .A2(g12382), .ZN(g21194) );
AND2_X4 U_g21195 ( .A1(g20212), .A2(g12385), .ZN(g21195) );
AND3_X4 U_I27761 ( .A1(g19411), .A2(g19382), .A3(g19352), .ZN(I27761) );
AND3_X4 U_g21196 ( .A1(g19329), .A2(g19313), .A3(I27761), .ZN(g21196) );
AND2_X4 U_g21197 ( .A1(g5912), .A2(g19330), .ZN(g21197) );
AND2_X4 U_g21198 ( .A1(g19534), .A2(g14601), .ZN(g21198) );
AND2_X4 U_g21203 ( .A1(g20178), .A2(g12409), .ZN(g21203) );
AND3_X4 U_I27772 ( .A1(g19314), .A2(g19501), .A3(g19480), .ZN(I27772) );
AND3_X4 U_g21207 ( .A1(g19456), .A2(g19430), .A3(I27772), .ZN(g21207) );
AND3_X4 U_g21208 ( .A1(g20150), .A2(g16619), .A3(g16586), .ZN(g21208) );
AND2_X4 U_g21209 ( .A1(g20273), .A2(g12412), .ZN(g21209) );
AND2_X4 U_g21210 ( .A1(g20242), .A2(g12415), .ZN(g21210) );
AND2_X4 U_g21218 ( .A1(g20212), .A2(g12421), .ZN(g21218) );
AND2_X4 U_g21226 ( .A1(g20242), .A2(g12426), .ZN(g21226) );
AND3_X4 U_g21229 ( .A1(g19578), .A2(g14797), .A3(g16665), .ZN(g21229) );
AND3_X4 U_g21234 ( .A1(g19608), .A2(g14849), .A3(g16686), .ZN(g21234) );
AND3_X4 U_g21243 ( .A1(g19641), .A2(g14922), .A3(g16712), .ZN(g21243) );
AND2_X4 U_g21245 ( .A1(g20299), .A2(g14837), .ZN(g21245) );
AND3_X4 U_g21251 ( .A1(g19681), .A2(g15003), .A3(g16743), .ZN(g21251) );
AND2_X4 U_g21252 ( .A1(g19578), .A2(g14895), .ZN(g21252) );
AND2_X4 U_g21254 ( .A1(g20318), .A2(g14910), .ZN(g21254) );
AND3_X4 U_g21259 ( .A1(g20299), .A2(g16722), .A3(g16682), .ZN(g21259) );
AND2_X4 U_g21260 ( .A1(g19608), .A2(g14976), .ZN(g21260) );
AND2_X4 U_g21262 ( .A1(g20337), .A2(g14991), .ZN(g21262) );
AND3_X4 U_g21267 ( .A1(g20318), .A2(g16764), .A3(g16708), .ZN(g21267) );
AND2_X4 U_g21268 ( .A1(g19641), .A2(g15065), .ZN(g21268) );
AND2_X4 U_g21270 ( .A1(g20357), .A2(g15080), .ZN(g21270) );
AND3_X4 U_g21276 ( .A1(g20337), .A2(g16791), .A3(g16739), .ZN(g21276) );
AND2_X4 U_g21277 ( .A1(g19681), .A2(g15161), .ZN(g21277) );
AND3_X4 U_g21283 ( .A1(g20357), .A2(g16820), .A3(g16781), .ZN(g21283) );
AND2_X4 U_g21284 ( .A1(g9356), .A2(g20269), .ZN(g21284) );
AND2_X4 U_g21290 ( .A1(g9356), .A2(g20278), .ZN(g21290) );
AND2_X4 U_g21291 ( .A1(g9293), .A2(g20279), .ZN(g21291) );
AND2_X4 U_g21292 ( .A1(g9453), .A2(g20281), .ZN(g21292) );
AND2_X4 U_g21298 ( .A1(g9356), .A2(g20286), .ZN(g21298) );
AND2_X4 U_g21299 ( .A1(g9293), .A2(g20287), .ZN(g21299) );
AND2_X4 U_g21300 ( .A1(g9232), .A2(g20288), .ZN(g21300) );
AND2_X4 U_g21301 ( .A1(g9453), .A2(g20289), .ZN(g21301) );
AND2_X4 U_g21302 ( .A1(g9374), .A2(g20290), .ZN(g21302) );
AND2_X4 U_g21303 ( .A1(g9595), .A2(g20292), .ZN(g21303) );
AND2_X4 U_g21304 ( .A1(g9293), .A2(g20296), .ZN(g21304) );
AND2_X4 U_g21305 ( .A1(g9232), .A2(g20297), .ZN(g21305) );
AND2_X4 U_g21306 ( .A1(g9187), .A2(g20298), .ZN(g21306) );
AND2_X4 U_g21307 ( .A1(g9453), .A2(g20302), .ZN(g21307) );
AND2_X4 U_g21308 ( .A1(g9374), .A2(g20303), .ZN(g21308) );
AND2_X4 U_g21309 ( .A1(g9310), .A2(g20304), .ZN(g21309) );
AND2_X4 U_g21310 ( .A1(g9595), .A2(g20305), .ZN(g21310) );
AND2_X4 U_g21311 ( .A1(g9471), .A2(g20306), .ZN(g21311) );
AND2_X4 U_g21312 ( .A1(g9737), .A2(g20308), .ZN(g21312) );
AND2_X4 U_g21313 ( .A1(g9232), .A2(g20311), .ZN(g21313) );
AND2_X4 U_g21314 ( .A1(g9187), .A2(g20312), .ZN(g21314) );
AND2_X4 U_g21315 ( .A1(g9161), .A2(g20313), .ZN(g21315) );
AND2_X4 U_g21319 ( .A1(g9374), .A2(g20315), .ZN(g21319) );
AND2_X4 U_g21320 ( .A1(g9310), .A2(g20316), .ZN(g21320) );
AND2_X4 U_g21321 ( .A1(g9248), .A2(g20317), .ZN(g21321) );
AND2_X4 U_g21322 ( .A1(g9595), .A2(g20321), .ZN(g21322) );
AND2_X4 U_g21323 ( .A1(g9471), .A2(g20322), .ZN(g21323) );
AND2_X4 U_g21324 ( .A1(g9391), .A2(g20323), .ZN(g21324) );
AND2_X4 U_g21325 ( .A1(g9737), .A2(g20324), .ZN(g21325) );
AND2_X4 U_g21326 ( .A1(g9613), .A2(g20325), .ZN(g21326) );
AND2_X4 U_g21328 ( .A1(g9187), .A2(g20327), .ZN(g21328) );
AND2_X4 U_g21329 ( .A1(g9161), .A2(g20328), .ZN(g21329) );
AND2_X4 U_g21330 ( .A1(g9150), .A2(g20329), .ZN(g21330) );
AND2_X4 U_g21334 ( .A1(g9310), .A2(g20330), .ZN(g21334) );
AND2_X4 U_g21335 ( .A1(g9248), .A2(g20331), .ZN(g21335) );
AND2_X4 U_g21336 ( .A1(g9203), .A2(g20332), .ZN(g21336) );
AND2_X4 U_g21337 ( .A1(g9471), .A2(g20334), .ZN(g21337) );
AND2_X4 U_g21338 ( .A1(g9391), .A2(g20335), .ZN(g21338) );
AND2_X4 U_g21339 ( .A1(g9326), .A2(g20336), .ZN(g21339) );
AND2_X4 U_g21340 ( .A1(g9737), .A2(g20340), .ZN(g21340) );
AND2_X4 U_g21341 ( .A1(g9613), .A2(g20341), .ZN(g21341) );
AND2_X4 U_g21342 ( .A1(g9488), .A2(g20342), .ZN(g21342) );
AND2_X4 U_g21343 ( .A1(g9161), .A2(g20344), .ZN(g21343) );
AND2_X4 U_g21344 ( .A1(g9150), .A2(g20345), .ZN(g21344) );
AND2_X4 U_g21345 ( .A1(g15096), .A2(g20346), .ZN(g21345) );
AND2_X4 U_g21349 ( .A1(g9248), .A2(g20347), .ZN(g21349) );
AND2_X4 U_g21350 ( .A1(g9203), .A2(g20348), .ZN(g21350) );
AND2_X4 U_g21351 ( .A1(g9174), .A2(g20349), .ZN(g21351) );
AND2_X4 U_g21352 ( .A1(g9391), .A2(g20350), .ZN(g21352) );
AND2_X4 U_g21353 ( .A1(g9326), .A2(g20351), .ZN(g21353) );
AND2_X4 U_g21354 ( .A1(g9264), .A2(g20352), .ZN(g21354) );
AND2_X4 U_g21355 ( .A1(g9613), .A2(g20354), .ZN(g21355) );
AND2_X4 U_g21356 ( .A1(g9488), .A2(g20355), .ZN(g21356) );
AND2_X4 U_g21357 ( .A1(g9407), .A2(g20356), .ZN(g21357) );
AND2_X4 U_g21360 ( .A1(g9507), .A2(g20361), .ZN(g21360) );
AND2_X4 U_g21361 ( .A1(g9150), .A2(g20362), .ZN(g21361) );
AND2_X4 U_g21362 ( .A1(g15096), .A2(g20363), .ZN(g21362) );
AND2_X4 U_g21363 ( .A1(g15022), .A2(g20364), .ZN(g21363) );
AND2_X4 U_g21367 ( .A1(g9203), .A2(g20366), .ZN(g21367) );
AND2_X4 U_g21368 ( .A1(g9174), .A2(g20367), .ZN(g21368) );
AND2_X4 U_g21369 ( .A1(g15188), .A2(g20368), .ZN(g21369) );
AND2_X4 U_g21370 ( .A1(g9326), .A2(g20369), .ZN(g21370) );
AND2_X4 U_g21371 ( .A1(g9264), .A2(g20370), .ZN(g21371) );
AND2_X4 U_g21372 ( .A1(g9216), .A2(g20371), .ZN(g21372) );
AND2_X4 U_g21373 ( .A1(g9488), .A2(g20372), .ZN(g21373) );
AND2_X4 U_g21374 ( .A1(g9407), .A2(g20373), .ZN(g21374) );
AND2_X4 U_g21375 ( .A1(g9342), .A2(g20374), .ZN(g21375) );
AND2_X4 U_g21378 ( .A1(g9507), .A2(g20378), .ZN(g21378) );
AND2_X4 U_g21379 ( .A1(g9427), .A2(g20379), .ZN(g21379) );
AND2_X4 U_g21380 ( .A1(g15096), .A2(g20380), .ZN(g21380) );
AND2_X4 U_g21381 ( .A1(g15022), .A2(g20381), .ZN(g21381) );
AND2_X4 U_g21388 ( .A1(g6201), .A2(g19657), .ZN(g21388) );
AND2_X4 U_g21389 ( .A1(g9649), .A2(g20384), .ZN(g21389) );
AND2_X4 U_g21390 ( .A1(g9174), .A2(g20385), .ZN(g21390) );
AND2_X4 U_g21391 ( .A1(g15188), .A2(g20386), .ZN(g21391) );
AND2_X4 U_g21392 ( .A1(g15118), .A2(g20387), .ZN(g21392) );
AND2_X4 U_g21393 ( .A1(g9264), .A2(g20389), .ZN(g21393) );
AND2_X4 U_g21394 ( .A1(g9216), .A2(g20390), .ZN(g21394) );
AND2_X4 U_g21395 ( .A1(g15274), .A2(g20391), .ZN(g21395) );
AND2_X4 U_g21396 ( .A1(g9407), .A2(g20392), .ZN(g21396) );
AND2_X4 U_g21397 ( .A1(g9342), .A2(g20393), .ZN(g21397) );
AND2_X4 U_g21398 ( .A1(g9277), .A2(g20394), .ZN(g21398) );
AND2_X4 U_g21401 ( .A1(g9507), .A2(g20397), .ZN(g21401) );
AND2_X4 U_g21402 ( .A1(g9427), .A2(g20398), .ZN(g21402) );
AND2_X4 U_g21403 ( .A1(g15022), .A2(g20399), .ZN(g21403) );
AND2_X4 U_g21410 ( .A1(g6363), .A2(g20402), .ZN(g21410) );
AND2_X4 U_g21411 ( .A1(g9649), .A2(g20403), .ZN(g21411) );
AND2_X4 U_g21412 ( .A1(g9569), .A2(g20404), .ZN(g21412) );
AND2_X4 U_g21413 ( .A1(g15188), .A2(g20405), .ZN(g21413) );
AND2_X4 U_g21414 ( .A1(g15118), .A2(g20406), .ZN(g21414) );
AND2_X4 U_g21418 ( .A1(g6290), .A2(g19705), .ZN(g21418) );
AND2_X4 U_g21419 ( .A1(g9795), .A2(g20409), .ZN(g21419) );
AND2_X4 U_g21420 ( .A1(g9216), .A2(g20410), .ZN(g21420) );
AND2_X4 U_g21421 ( .A1(g15274), .A2(g20411), .ZN(g21421) );
AND2_X4 U_g21422 ( .A1(g15210), .A2(g20412), .ZN(g21422) );
AND2_X4 U_g21423 ( .A1(g9342), .A2(g20414), .ZN(g21423) );
AND2_X4 U_g21424 ( .A1(g9277), .A2(g20415), .ZN(g21424) );
AND2_X4 U_g21425 ( .A1(g15366), .A2(g20416), .ZN(g21425) );
AND2_X4 U_g21428 ( .A1(g9427), .A2(g20420), .ZN(g21428) );
AND2_X4 U_g21438 ( .A1(g9649), .A2(g20422), .ZN(g21438) );
AND2_X4 U_g21439 ( .A1(g9569), .A2(g20423), .ZN(g21439) );
AND2_X4 U_g21440 ( .A1(g15118), .A2(g20424), .ZN(g21440) );
AND2_X4 U_g21444 ( .A1(g6568), .A2(g20427), .ZN(g21444) );
AND2_X4 U_g21445 ( .A1(g9795), .A2(g20428), .ZN(g21445) );
AND2_X4 U_g21446 ( .A1(g9711), .A2(g20429), .ZN(g21446) );
AND2_X4 U_g21447 ( .A1(g15274), .A2(g20430), .ZN(g21447) );
AND2_X4 U_g21448 ( .A1(g15210), .A2(g20431), .ZN(g21448) );
AND2_X4 U_g21452 ( .A1(g6427), .A2(g19749), .ZN(g21452) );
AND2_X4 U_g21453 ( .A1(g9941), .A2(g20434), .ZN(g21453) );
AND2_X4 U_g21454 ( .A1(g9277), .A2(g20435), .ZN(g21454) );
AND2_X4 U_g21455 ( .A1(g15366), .A2(g20436), .ZN(g21455) );
AND2_X4 U_g21456 ( .A1(g15296), .A2(g20437), .ZN(g21456) );
AND2_X4 U_g21476 ( .A1(g9569), .A2(g20442), .ZN(g21476) );
AND2_X4 U_g21480 ( .A1(g9795), .A2(g20444), .ZN(g21480) );
AND2_X4 U_g21481 ( .A1(g9711), .A2(g20445), .ZN(g21481) );
AND2_X4 U_g21482 ( .A1(g15210), .A2(g20446), .ZN(g21482) );
AND2_X4 U_g21486 ( .A1(g6832), .A2(g20449), .ZN(g21486) );
AND2_X4 U_g21487 ( .A1(g9941), .A2(g20450), .ZN(g21487) );
AND2_X4 U_g21488 ( .A1(g9857), .A2(g20451), .ZN(g21488) );
AND2_X4 U_g21489 ( .A1(g15366), .A2(g20452), .ZN(g21489) );
AND2_X4 U_g21490 ( .A1(g15296), .A2(g20453), .ZN(g21490) );
AND2_X4 U_g21494 ( .A1(g6632), .A2(g19792), .ZN(g21494) );
AND2_X4 U_g21497 ( .A1(g3006), .A2(g20456), .ZN(g21497) );
AND2_X4 U_g21517 ( .A1(g9711), .A2(g20461), .ZN(g21517) );
AND2_X4 U_g21521 ( .A1(g9941), .A2(g20463), .ZN(g21521) );
AND2_X4 U_g21522 ( .A1(g9857), .A2(g20464), .ZN(g21522) );
AND2_X4 U_g21523 ( .A1(g15296), .A2(g20465), .ZN(g21523) );
AND2_X4 U_g21527 ( .A1(g7134), .A2(g20468), .ZN(g21527) );
AND3_X4 U_I28068 ( .A1(g17802), .A2(g18265), .A3(g17882), .ZN(I28068) );
AND4_X4 U_g21533 ( .A1(g17724), .A2(g18179), .A3(g19799), .A4(I28068), .ZN(g21533) );
AND2_X4 U_g21553 ( .A1(g9857), .A2(g20476), .ZN(g21553) );
AND3_X4 U_I28096 ( .A1(g13907), .A2(g14238), .A3(g13946), .ZN(I28096) );
AND4_X4 U_g21564 ( .A1(g13886), .A2(g14153), .A3(g19799), .A4(I28096), .ZN(g21564) );
AND3_X4 U_I28103 ( .A1(g17914), .A2(g18358), .A3(g17993), .ZN(I28103) );
AND4_X4 U_g21569 ( .A1(g17825), .A2(g18286), .A3(g19843), .A4(I28103), .ZN(g21569) );
AND2_X4 U_g21589 ( .A1(g3002), .A2(g19890), .ZN(g21589) );
AND3_X4 U_g21593 ( .A1(g16498), .A2(g19484), .A3(g14071), .ZN(g21593) );
AND3_X4 U_I28126 ( .A1(g13963), .A2(g14360), .A3(g14016), .ZN(I28126) );
AND4_X4 U_g21597 ( .A1(g13927), .A2(g14268), .A3(g19843), .A4(I28126), .ZN(g21597) );
AND3_X4 U_I28133 ( .A1(g18025), .A2(g18453), .A3(g18110), .ZN(I28133) );
AND4_X4 U_g21602 ( .A1(g17937), .A2(g18379), .A3(g19876), .A4(I28133), .ZN(g21602) );
AND2_X4 U_g21610 ( .A1(g7522), .A2(g20490), .ZN(g21610) );
AND2_X4 U_g21611 ( .A1(g7471), .A2(g19915), .ZN(g21611) );
AND3_X4 U_g21622 ( .A1(g16520), .A2(g19505), .A3(g14186), .ZN(g21622) );
AND3_X4 U_I28155 ( .A1(g14033), .A2(g14472), .A3(g14107), .ZN(I28155) );
AND4_X4 U_g21626 ( .A1(g13983), .A2(g14390), .A3(g19876), .A4(I28155), .ZN(g21626) );
AND3_X4 U_I28162 ( .A1(g18142), .A2(g18526), .A3(g18226), .ZN(I28162) );
AND4_X4 U_g21631 ( .A1(g18048), .A2(g18474), .A3(g19907), .A4(I28162), .ZN(g21631) );
AND2_X4 U_g21635 ( .A1(g7549), .A2(g20496), .ZN(g21635) );
AND2_X4 U_g21639 ( .A1(g3398), .A2(g20500), .ZN(g21639) );
AND3_X4 U_g21650 ( .A1(g16551), .A2(g19524), .A3(g14301), .ZN(g21650) );
AND3_X4 U_I28181 ( .A1(g14124), .A2(g14559), .A3(g14222), .ZN(I28181) );
AND4_X4 U_g21654 ( .A1(g14053), .A2(g14502), .A3(g19907), .A4(I28181), .ZN(g21654) );
AND2_X4 U_g21658 ( .A1(g2896), .A2(g20501), .ZN(g21658) );
AND2_X4 U_g21666 ( .A1(g3398), .A2(g20504), .ZN(g21666) );
AND2_X4 U_g21670 ( .A1(g3554), .A2(g20505), .ZN(g21670) );
AND3_X4 U_g21681 ( .A1(g16583), .A2(g19534), .A3(g14423), .ZN(g21681) );
AND2_X4 U_g21687 ( .A1(g3398), .A2(g20516), .ZN(g21687) );
AND2_X4 U_g21695 ( .A1(g3554), .A2(g20517), .ZN(g21695) );
AND2_X4 U_g21699 ( .A1(g3710), .A2(g20518), .ZN(g21699) );
AND2_X4 U_g21707 ( .A1(g2892), .A2(g19978), .ZN(g21707) );
AND2_X4 U_g21723 ( .A1(g3554), .A2(g20534), .ZN(g21723) );
AND2_X4 U_g21731 ( .A1(g3710), .A2(g20535), .ZN(g21731) );
AND2_X4 U_g21735 ( .A1(g3866), .A2(g20536), .ZN(g21735) );
AND2_X4 U_g21749 ( .A1(g3710), .A2(g20553), .ZN(g21749) );
AND2_X4 U_g21757 ( .A1(g3866), .A2(g20554), .ZN(g21757) );
AND2_X4 U_g21758 ( .A1(g7607), .A2(g20045), .ZN(g21758) );
AND2_X4 U_g21773 ( .A1(g3866), .A2(g19078), .ZN(g21773) );
AND3_X4 U_g21805 ( .A1(g16679), .A2(g19578), .A3(g14776), .ZN(g21805) );
AND3_X4 U_g21812 ( .A1(g16705), .A2(g19608), .A3(g14811), .ZN(g21812) );
AND3_X4 U_g21818 ( .A1(g16736), .A2(g19641), .A3(g14863), .ZN(g21818) );
AND3_X4 U_g21822 ( .A1(g16778), .A2(g19681), .A3(g14936), .ZN(g21822) );
AND2_X4 U_g21891 ( .A1(g19302), .A2(g11749), .ZN(g21891) );
AND2_X4 U_g21892 ( .A1(g19288), .A2(g13011), .ZN(g21892) );
AND2_X4 U_g21899 ( .A1(g19323), .A2(g11749), .ZN(g21899) );
AND2_X4 U_g21900 ( .A1(g19306), .A2(g13011), .ZN(g21900) );
AND2_X4 U_g21906 ( .A1(g5715), .A2(g20513), .ZN(g21906) );
AND2_X4 U_g21911 ( .A1(g19350), .A2(g11749), .ZN(g21911) );
AND2_X4 U_g21912 ( .A1(g19327), .A2(g13011), .ZN(g21912) );
AND2_X4 U_g21913 ( .A1(g4456), .A2(g20519), .ZN(g21913) );
AND2_X4 U_g21920 ( .A1(g5773), .A2(g20531), .ZN(g21920) );
AND2_X4 U_g21925 ( .A1(g19384), .A2(g11749), .ZN(g21925) );
AND2_X4 U_g21926 ( .A1(g19354), .A2(g13011), .ZN(g21926) );
AND2_X4 U_g21931 ( .A1(g4632), .A2(g20539), .ZN(g21931) );
AND2_X4 U_g21938 ( .A1(g5832), .A2(g20550), .ZN(g21938) );
AND2_X4 U_g21990 ( .A1(g291), .A2(g21187), .ZN(g21990) );
AND2_X4 U_g22004 ( .A1(g978), .A2(g21202), .ZN(g22004) );
AND2_X4 U_g22015 ( .A1(g1672), .A2(g21217), .ZN(g22015) );
AND2_X4 U_g22020 ( .A1(g2366), .A2(g21225), .ZN(g22020) );
AND3_X4 U_I28582 ( .A1(g19141), .A2(g21133), .A3(g21116), .ZN(I28582) );
AND4_X4 U_g22036 ( .A1(g21104), .A2(g21095), .A3(g21084), .A4(I28582), .ZN(g22036) );
AND3_X4 U_I28594 ( .A1(g21167), .A2(g21147), .A3(g21134), .ZN(I28594) );
AND4_X4 U_g22046 ( .A1(g21117), .A2(g21105), .A3(g21096), .A4(I28594), .ZN(g22046) );
AND3_X4 U_I28609 ( .A1(g21183), .A2(g21168), .A3(g21148), .ZN(I28609) );
AND4_X4 U_g22062 ( .A1(g21135), .A2(g21118), .A3(g21106), .A4(I28609), .ZN(g22062) );
AND2_X4 U_g22187 ( .A1(g21564), .A2(g20986), .ZN(g22187) );
AND2_X4 U_g22196 ( .A1(g21597), .A2(g21012), .ZN(g22196) );
AND2_X4 U_g22201 ( .A1(g21271), .A2(g16881), .ZN(g22201) );
AND2_X4 U_g22202 ( .A1(g21626), .A2(g21036), .ZN(g22202) );
AND2_X4 U_g22206 ( .A1(g21895), .A2(g11976), .ZN(g22206) );
AND2_X4 U_g22207 ( .A1(g21278), .A2(g16910), .ZN(g22207) );
AND2_X4 U_g22208 ( .A1(g21654), .A2(g21057), .ZN(g22208) );
AND2_X4 U_g22211 ( .A1(g21661), .A2(g12027), .ZN(g22211) );
AND2_X4 U_g22214 ( .A1(g21907), .A2(g12045), .ZN(g22214) );
AND2_X4 U_g22215 ( .A1(g21285), .A2(g16940), .ZN(g22215) );
AND2_X4 U_g22220 ( .A1(g21690), .A2(g12091), .ZN(g22220) );
AND2_X4 U_g22223 ( .A1(g21921), .A2(g12109), .ZN(g22223) );
AND2_X4 U_g22224 ( .A1(g21293), .A2(g16971), .ZN(g22224) );
AND2_X4 U_g22228 ( .A1(g21716), .A2(g12136), .ZN(g22228) );
AND2_X4 U_g22229 ( .A1(g21661), .A2(g12139), .ZN(g22229) );
AND2_X4 U_g22235 ( .A1(g21726), .A2(g12163), .ZN(g22235) );
AND2_X4 U_g22238 ( .A1(g21939), .A2(g12181), .ZN(g22238) );
AND2_X4 U_g22244 ( .A1(g21742), .A2(g12198), .ZN(g22244) );
AND2_X4 U_g22245 ( .A1(g21690), .A2(g12201), .ZN(g22245) );
AND2_X4 U_g22250 ( .A1(g21752), .A2(g12225), .ZN(g22250) );
AND2_X4 U_g22254 ( .A1(g21716), .A2(g12239), .ZN(g22254) );
AND2_X4 U_g22255 ( .A1(g21661), .A2(g12242), .ZN(g22255) );
AND2_X4 U_g22264 ( .A1(g21766), .A2(g12253), .ZN(g22264) );
AND2_X4 U_g22265 ( .A1(g21726), .A2(g12256), .ZN(g22265) );
AND2_X4 U_g22270 ( .A1(g92), .A2(g21529), .ZN(g22270) );
AND2_X4 U_g22272 ( .A1(g21742), .A2(g12282), .ZN(g22272) );
AND2_X4 U_g22273 ( .A1(g21690), .A2(g12285), .ZN(g22273) );
AND2_X4 U_g22281 ( .A1(g21782), .A2(g12296), .ZN(g22281) );
AND2_X4 U_g22282 ( .A1(g21752), .A2(g12299), .ZN(g22282) );
AND2_X4 U_g22285 ( .A1(g21716), .A2(g12312), .ZN(g22285) );
AND2_X4 U_g22289 ( .A1(g780), .A2(g21565), .ZN(g22289) );
AND2_X4 U_g22291 ( .A1(g21766), .A2(g12318), .ZN(g22291) );
AND2_X4 U_g22292 ( .A1(g21726), .A2(g12321), .ZN(g22292) );
AND2_X4 U_g22305 ( .A1(g21742), .A2(g12340), .ZN(g22305) );
AND2_X4 U_g22309 ( .A1(g1466), .A2(g21598), .ZN(g22309) );
AND2_X4 U_g22311 ( .A1(g21782), .A2(g12346), .ZN(g22311) );
AND2_X4 U_g22312 ( .A1(g21752), .A2(g12349), .ZN(g22312) );
AND2_X4 U_g22333 ( .A1(g21766), .A2(g12370), .ZN(g22333) );
AND2_X4 U_g22337 ( .A1(g2160), .A2(g21627), .ZN(g22337) );
AND2_X4 U_g22340 ( .A1(g88), .A2(g21184), .ZN(g22340) );
AND2_X4 U_g22358 ( .A1(g21782), .A2(g12389), .ZN(g22358) );
AND2_X4 U_g22363 ( .A1(g776), .A2(g21199), .ZN(g22363) );
AND2_X4 U_g22383 ( .A1(g1462), .A2(g21214), .ZN(g22383) );
AND2_X4 U_g22398 ( .A1(g2156), .A2(g21222), .ZN(g22398) );
AND2_X4 U_g22483 ( .A1(g646), .A2(g21861), .ZN(g22483) );
AND2_X4 U_g22515 ( .A1(g13873), .A2(g21382), .ZN(g22515) );
AND2_X4 U_g22516 ( .A1(g20885), .A2(g17442), .ZN(g22516) );
AND2_X4 U_g22517 ( .A1(g21895), .A2(g12608), .ZN(g22517) );
AND2_X4 U_g22526 ( .A1(g1332), .A2(g21867), .ZN(g22526) );
AND2_X4 U_g22546 ( .A1(g13886), .A2(g21404), .ZN(g22546) );
AND2_X4 U_g22555 ( .A1(g13895), .A2(g21415), .ZN(g22555) );
AND2_X4 U_g22556 ( .A1(g20904), .A2(g17523), .ZN(g22556) );
AND2_X4 U_g22557 ( .A1(g21907), .A2(g12654), .ZN(g22557) );
AND2_X4 U_g22566 ( .A1(g2026), .A2(g21872), .ZN(g22566) );
AND2_X4 U_g22577 ( .A1(g13907), .A2(g21429), .ZN(g22577) );
AND2_X4 U_g22581 ( .A1(g21895), .A2(g12699), .ZN(g22581) );
AND2_X4 U_g22587 ( .A1(g13927), .A2(g21441), .ZN(g22587) );
AND2_X4 U_g22595 ( .A1(g13936), .A2(g21449), .ZN(g22595) );
AND2_X4 U_g22596 ( .A1(g20928), .A2(g17613), .ZN(g22596) );
AND2_X4 U_g22597 ( .A1(g21921), .A2(g12708), .ZN(g22597) );
AND2_X4 U_g22606 ( .A1(g2720), .A2(g21876), .ZN(g22606) );
AND2_X4 U_g22607 ( .A1(g13946), .A2(g21458), .ZN(g22607) );
AND2_X4 U_g22610 ( .A1(g660), .A2(g21473), .ZN(g22610) );
AND2_X4 U_g22614 ( .A1(g13963), .A2(g21477), .ZN(g22614) );
AND2_X4 U_g22618 ( .A1(g21907), .A2(g12756), .ZN(g22618) );
AND2_X4 U_g22624 ( .A1(g13983), .A2(g21483), .ZN(g22624) );
AND2_X4 U_g22632 ( .A1(g13992), .A2(g21491), .ZN(g22632) );
AND2_X4 U_g22633 ( .A1(g20956), .A2(g17710), .ZN(g22633) );
AND2_X4 U_g22634 ( .A1(g21939), .A2(g12765), .ZN(g22634) );
AND2_X4 U_g22637 ( .A1(g20841), .A2(g10927), .ZN(g22637) );
AND2_X4 U_g22638 ( .A1(g14001), .A2(g21498), .ZN(g22638) );
AND2_X4 U_g22643 ( .A1(g14016), .A2(g21505), .ZN(g22643) );
AND2_X4 U_g22646 ( .A1(g1346), .A2(g21514), .ZN(g22646) );
AND2_X4 U_g22650 ( .A1(g14033), .A2(g21518), .ZN(g22650) );
AND2_X4 U_g22654 ( .A1(g21921), .A2(g12798), .ZN(g22654) );
AND2_X4 U_g22660 ( .A1(g14053), .A2(g21524), .ZN(g22660) );
AND2_X4 U_g22665 ( .A1(g20920), .A2(g6153), .ZN(g22665) );
AND2_X4 U_g22666 ( .A1(g21825), .A2(g20014), .ZN(g22666) );
AND2_X4 U_g22667 ( .A1(g14062), .A2(g21530), .ZN(g22667) );
AND2_X4 U_g22674 ( .A1(g14092), .A2(g21537), .ZN(g22674) );
AND2_X4 U_g22679 ( .A1(g14107), .A2(g21541), .ZN(g22679) );
AND2_X4 U_g22682 ( .A1(g2040), .A2(g21550), .ZN(g22682) );
AND2_X4 U_g22686 ( .A1(g14124), .A2(g21554), .ZN(g22686) );
AND2_X4 U_g22690 ( .A1(g21939), .A2(g12837), .ZN(g22690) );
AND2_X4 U_g22699 ( .A1(g7338), .A2(g21883), .ZN(g22699) );
AND2_X4 U_g22700 ( .A1(g7146), .A2(g21558), .ZN(g22700) );
AND2_X4 U_g22701 ( .A1(g18174), .A2(g21561), .ZN(g22701) );
AND2_X4 U_g22707 ( .A1(g14177), .A2(g21566), .ZN(g22707) );
AND2_X4 U_g22714 ( .A1(g14207), .A2(g21573), .ZN(g22714) );
AND2_X4 U_g22719 ( .A1(g14222), .A2(g21577), .ZN(g22719) );
AND2_X4 U_g22722 ( .A1(g2734), .A2(g21586), .ZN(g22722) );
AND2_X4 U_g22726 ( .A1(g3036), .A2(g21886), .ZN(g22726) );
AND2_X4 U_g22727 ( .A1(g14238), .A2(g21590), .ZN(g22727) );
AND2_X4 U_g22732 ( .A1(g18281), .A2(g21594), .ZN(g22732) );
AND2_X4 U_g22738 ( .A1(g14292), .A2(g21599), .ZN(g22738) );
AND2_X4 U_g22745 ( .A1(g14322), .A2(g21606), .ZN(g22745) );
AND2_X4 U_g22754 ( .A1(g14342), .A2(g21612), .ZN(g22754) );
AND2_X4 U_g22759 ( .A1(g14360), .A2(g21619), .ZN(g22759) );
AND2_X4 U_g22764 ( .A1(g18374), .A2(g21623), .ZN(g22764) );
AND2_X4 U_g22770 ( .A1(g14414), .A2(g21628), .ZN(g22770) );
AND2_X4 U_g22788 ( .A1(g14454), .A2(g21640), .ZN(g22788) );
AND2_X4 U_g22793 ( .A1(g14472), .A2(g21647), .ZN(g22793) );
AND2_X4 U_g22798 ( .A1(g18469), .A2(g21651), .ZN(g22798) );
AND2_X4 U_g22804 ( .A1(g2920), .A2(g21655), .ZN(g22804) );
AND2_X4 U_g22830 ( .A1(g14541), .A2(g21671), .ZN(g22830) );
AND2_X4 U_g22835 ( .A1(g14559), .A2(g21678), .ZN(g22835) );
AND2_X4 U_g22841 ( .A1(g7583), .A2(g21902), .ZN(g22841) );
AND2_X4 U_g22842 ( .A1(g3032), .A2(g21682), .ZN(g22842) );
AND2_X4 U_g22869 ( .A1(g14596), .A2(g21700), .ZN(g22869) );
AND2_X4 U_g22874 ( .A1(g7587), .A2(g21708), .ZN(g22874) );
AND2_X4 U_g22906 ( .A1(g2924), .A2(g21927), .ZN(g22906) );
AND2_X4 U_g22984 ( .A1(g16840), .A2(g21400), .ZN(g22984) );
AND2_X4 U_g23104 ( .A1(g20842), .A2(g15859), .ZN(g23104) );
AND2_X4 U_g23106 ( .A1(g5857), .A2(g21050), .ZN(g23106) );
AND2_X4 U_g23118 ( .A1(g20850), .A2(g15890), .ZN(g23118) );
AND2_X4 U_g23119 ( .A1(g5904), .A2(g21069), .ZN(g23119) );
AND2_X4 U_g23127 ( .A1(g20858), .A2(g15923), .ZN(g23127) );
AND2_X4 U_g23128 ( .A1(g5943), .A2(g21079), .ZN(g23128) );
AND2_X4 U_g23138 ( .A1(g20866), .A2(g15952), .ZN(g23138) );
AND2_X4 U_g23139 ( .A1(g5977), .A2(g21093), .ZN(g23139) );
AND2_X4 U_g23409 ( .A1(g21533), .A2(g22408), .ZN(g23409) );
AND2_X4 U_g23414 ( .A1(g21569), .A2(g22421), .ZN(g23414) );
AND2_X4 U_g23419 ( .A1(g22755), .A2(g19577), .ZN(g23419) );
AND2_X4 U_g23423 ( .A1(g21602), .A2(g22443), .ZN(g23423) );
AND2_X4 U_g23428 ( .A1(g22789), .A2(g19607), .ZN(g23428) );
AND2_X4 U_g23432 ( .A1(g21631), .A2(g22476), .ZN(g23432) );
AND2_X4 U_g23434 ( .A1(g22831), .A2(g19640), .ZN(g23434) );
AND2_X4 U_g23440 ( .A1(g22870), .A2(g19680), .ZN(g23440) );
AND2_X4 U_g23451 ( .A1(g18552), .A2(g22547), .ZN(g23451) );
AND2_X4 U_g23458 ( .A1(g18602), .A2(g22588), .ZN(g23458) );
AND2_X4 U_g23462 ( .A1(g17988), .A2(g22609), .ZN(g23462) );
AND2_X4 U_g23467 ( .A1(g18634), .A2(g22625), .ZN(g23467) );
AND2_X4 U_g23471 ( .A1(g18105), .A2(g22645), .ZN(g23471) );
AND2_X4 U_g23476 ( .A1(g18643), .A2(g22661), .ZN(g23476) );
AND2_X4 U_g23483 ( .A1(g22945), .A2(g8847), .ZN(g23483) );
AND2_X4 U_g23484 ( .A1(g18221), .A2(g22681), .ZN(g23484) );
AND2_X4 U_g23494 ( .A1(g18328), .A2(g22721), .ZN(g23494) );
AND2_X4 U_g23496 ( .A1(g5802), .A2(g22300), .ZN(g23496) );
AND2_X4 U_g23510 ( .A1(g5890), .A2(g22753), .ZN(g23510) );
AND2_X4 U_g23512 ( .A1(g5858), .A2(g22328), .ZN(g23512) );
AND2_X4 U_g23525 ( .A1(g5929), .A2(g22787), .ZN(g23525) );
AND2_X4 U_g23527 ( .A1(g5905), .A2(g22353), .ZN(g23527) );
AND2_X4 U_g23536 ( .A1(g5963), .A2(g22829), .ZN(g23536) );
AND2_X4 U_g23538 ( .A1(g5944), .A2(g22376), .ZN(g23538) );
AND2_X4 U_g23544 ( .A1(g5992), .A2(g22868), .ZN(g23544) );
AND2_X4 U_g23547 ( .A1(g8062), .A2(g22405), .ZN(g23547) );
AND2_X4 U_g23550 ( .A1(g8132), .A2(g22409), .ZN(g23550) );
AND2_X4 U_g23551 ( .A1(g8135), .A2(g22412), .ZN(g23551) );
AND2_X4 U_g23552 ( .A1(g6136), .A2(g22415), .ZN(g23552) );
AND2_X4 U_g23554 ( .A1(g8147), .A2(g22418), .ZN(g23554) );
AND2_X4 U_g23558 ( .A1(g8200), .A2(g22422), .ZN(g23558) );
AND2_X4 U_g23559 ( .A1(g8203), .A2(g22425), .ZN(g23559) );
AND2_X4 U_g23560 ( .A1(g8206), .A2(g22428), .ZN(g23560) );
AND2_X4 U_g23563 ( .A1(g8218), .A2(g22431), .ZN(g23563) );
AND2_X4 U_g23564 ( .A1(g8221), .A2(g22434), .ZN(g23564) );
AND2_X4 U_g23565 ( .A1(g6146), .A2(g22437), .ZN(g23565) );
AND2_X4 U_g23567 ( .A1(g8233), .A2(g22440), .ZN(g23567) );
AND2_X4 U_g23571 ( .A1(g3931), .A2(g22445), .ZN(g23571) );
AND2_X4 U_g23572 ( .A1(g3934), .A2(g22448), .ZN(g23572) );
AND2_X4 U_g23573 ( .A1(g3937), .A2(g22451), .ZN(g23573) );
AND2_X4 U_g23577 ( .A1(g3957), .A2(g22455), .ZN(g23577) );
AND2_X4 U_g23578 ( .A1(g3960), .A2(g22458), .ZN(g23578) );
AND2_X4 U_g23579 ( .A1(g3963), .A2(g22461), .ZN(g23579) );
AND2_X4 U_g23582 ( .A1(g3975), .A2(g22464), .ZN(g23582) );
AND2_X4 U_g23583 ( .A1(g3978), .A2(g22467), .ZN(g23583) );
AND2_X4 U_g23584 ( .A1(g6167), .A2(g22470), .ZN(g23584) );
AND2_X4 U_g23586 ( .A1(g3990), .A2(g22473), .ZN(g23586) );
AND2_X4 U_g23590 ( .A1(g4009), .A2(g22477), .ZN(g23590) );
AND2_X4 U_g23591 ( .A1(g4012), .A2(g22480), .ZN(g23591) );
AND2_X4 U_g23592 ( .A1(g17640), .A2(g22986), .ZN(g23592) );
AND2_X4 U_g23593 ( .A1(g22845), .A2(g20365), .ZN(g23593) );
AND2_X4 U_g23598 ( .A1(g4038), .A2(g22484), .ZN(g23598) );
AND2_X4 U_g23599 ( .A1(g4041), .A2(g22487), .ZN(g23599) );
AND2_X4 U_g23600 ( .A1(g4044), .A2(g22490), .ZN(g23600) );
AND2_X4 U_g23604 ( .A1(g4064), .A2(g22494), .ZN(g23604) );
AND2_X4 U_g23605 ( .A1(g4067), .A2(g22497), .ZN(g23605) );
AND2_X4 U_g23606 ( .A1(g4070), .A2(g22500), .ZN(g23606) );
AND2_X4 U_g23609 ( .A1(g4082), .A2(g22503), .ZN(g23609) );
AND2_X4 U_g23610 ( .A1(g4085), .A2(g22506), .ZN(g23610) );
AND2_X4 U_g23611 ( .A1(g6194), .A2(g22509), .ZN(g23611) );
AND2_X4 U_g23615 ( .A1(g4107), .A2(g22512), .ZN(g23615) );
AND2_X4 U_g23616 ( .A1(g17724), .A2(g22988), .ZN(g23616) );
AND2_X4 U_g23617 ( .A1(g22810), .A2(g20382), .ZN(g23617) );
AND2_X4 U_g23618 ( .A1(g22608), .A2(g20383), .ZN(g23618) );
AND2_X4 U_g23622 ( .A1(g4136), .A2(g22520), .ZN(g23622) );
AND2_X4 U_g23623 ( .A1(g4139), .A2(g22523), .ZN(g23623) );
AND2_X4 U_g23624 ( .A1(g17741), .A2(g22989), .ZN(g23624) );
AND2_X4 U_g23625 ( .A1(g22880), .A2(g20388), .ZN(g23625) );
AND2_X4 U_g23630 ( .A1(g4165), .A2(g22527), .ZN(g23630) );
AND2_X4 U_g23631 ( .A1(g4168), .A2(g22530), .ZN(g23631) );
AND2_X4 U_g23632 ( .A1(g4171), .A2(g22533), .ZN(g23632) );
AND2_X4 U_g23636 ( .A1(g4191), .A2(g22537), .ZN(g23636) );
AND2_X4 U_g23637 ( .A1(g4194), .A2(g22540), .ZN(g23637) );
AND2_X4 U_g23638 ( .A1(g4197), .A2(g22543), .ZN(g23638) );
AND2_X4 U_g23639 ( .A1(g21825), .A2(g22805), .ZN(g23639) );
AND2_X4 U_g23643 ( .A1(g17802), .A2(g22991), .ZN(g23643) );
AND2_X4 U_g23659 ( .A1(g22784), .A2(g17500), .ZN(g23659) );
AND2_X4 U_g23664 ( .A1(g4246), .A2(g22552), .ZN(g23664) );
AND2_X4 U_g23665 ( .A1(g17825), .A2(g22995), .ZN(g23665) );
AND2_X4 U_g23666 ( .A1(g22851), .A2(g20407), .ZN(g23666) );
AND2_X4 U_g23667 ( .A1(g22644), .A2(g20408), .ZN(g23667) );
AND2_X4 U_g23671 ( .A1(g4275), .A2(g22560), .ZN(g23671) );
AND2_X4 U_g23672 ( .A1(g4278), .A2(g22563), .ZN(g23672) );
AND2_X4 U_g23673 ( .A1(g17842), .A2(g22996), .ZN(g23673) );
AND2_X4 U_g23674 ( .A1(g22915), .A2(g20413), .ZN(g23674) );
AND2_X4 U_g23679 ( .A1(g4304), .A2(g22567), .ZN(g23679) );
AND2_X4 U_g23680 ( .A1(g4307), .A2(g22570), .ZN(g23680) );
AND2_X4 U_g23681 ( .A1(g4310), .A2(g22573), .ZN(g23681) );
AND2_X4 U_g23686 ( .A1(g17882), .A2(g22998), .ZN(g23686) );
AND2_X4 U_g23687 ( .A1(g22668), .A2(g17570), .ZN(g23687) );
AND2_X4 U_g23689 ( .A1(g6513), .A2(g23001), .ZN(g23689) );
AND2_X4 U_g23693 ( .A1(g17914), .A2(g23002), .ZN(g23693) );
AND2_X4 U_g23709 ( .A1(g22826), .A2(g17591), .ZN(g23709) );
AND2_X4 U_g23714 ( .A1(g4401), .A2(g22592), .ZN(g23714) );
AND2_X4 U_g23715 ( .A1(g17937), .A2(g23006), .ZN(g23715) );
AND2_X4 U_g23716 ( .A1(g22886), .A2(g20432), .ZN(g23716) );
AND2_X4 U_g23717 ( .A1(g22680), .A2(g20433), .ZN(g23717) );
AND2_X4 U_g23721 ( .A1(g4430), .A2(g22600), .ZN(g23721) );
AND2_X4 U_g23722 ( .A1(g4433), .A2(g22603), .ZN(g23722) );
AND2_X4 U_g23723 ( .A1(g17954), .A2(g23007), .ZN(g23723) );
AND2_X4 U_g23724 ( .A1(g22940), .A2(g20438), .ZN(g23724) );
AND2_X4 U_g23726 ( .A1(g21825), .A2(g22843), .ZN(g23726) );
AND2_X4 U_g23734 ( .A1(g17974), .A2(g23008), .ZN(g23734) );
AND2_X4 U_g23735 ( .A1(g22949), .A2(g9450), .ZN(g23735) );
AND2_X4 U_g23740 ( .A1(g17993), .A2(g23012), .ZN(g23740) );
AND2_X4 U_g23741 ( .A1(g22708), .A2(g17667), .ZN(g23741) );
AND2_X4 U_g23743 ( .A1(g6777), .A2(g23015), .ZN(g23743) );
AND2_X4 U_g23747 ( .A1(g18025), .A2(g23016), .ZN(g23747) );
AND2_X4 U_g23763 ( .A1(g22865), .A2(g17688), .ZN(g23763) );
AND2_X4 U_g23768 ( .A1(g4570), .A2(g22629), .ZN(g23768) );
AND2_X4 U_g23769 ( .A1(g18048), .A2(g23020), .ZN(g23769) );
AND2_X4 U_g23770 ( .A1(g22921), .A2(g20454), .ZN(g23770) );
AND2_X4 U_g23771 ( .A1(g22720), .A2(g20455), .ZN(g23771) );
AND2_X4 U_g23772 ( .A1(g21825), .A2(g22875), .ZN(g23772) );
AND2_X4 U_g23776 ( .A1(g18074), .A2(g23021), .ZN(g23776) );
AND2_X4 U_g23777 ( .A1(g22949), .A2(g9528), .ZN(g23777) );
AND2_X4 U_g23778 ( .A1(g22954), .A2(g9531), .ZN(g23778) );
AND2_X4 U_g23789 ( .A1(g18091), .A2(g23024), .ZN(g23789) );
AND2_X4 U_g23790 ( .A1(g22958), .A2(g9592), .ZN(g23790) );
AND2_X4 U_g23795 ( .A1(g18110), .A2(g23028), .ZN(g23795) );
AND2_X4 U_g23796 ( .A1(g22739), .A2(g17767), .ZN(g23796) );
AND2_X4 U_g23798 ( .A1(g7079), .A2(g23031), .ZN(g23798) );
AND2_X4 U_g23802 ( .A1(g18142), .A2(g23032), .ZN(g23802) );
AND2_X4 U_g23818 ( .A1(g22900), .A2(g17788), .ZN(g23818) );
AND2_X4 U_g23820 ( .A1(g3013), .A2(g23036), .ZN(g23820) );
AND2_X4 U_g23822 ( .A1(g14148), .A2(g23037), .ZN(g23822) );
AND2_X4 U_g23824 ( .A1(g22949), .A2(g9641), .ZN(g23824) );
AND2_X4 U_g23825 ( .A1(g22954), .A2(g9644), .ZN(g23825) );
AND2_X4 U_g23829 ( .A1(g18190), .A2(g23038), .ZN(g23829) );
AND2_X4 U_g23830 ( .A1(g22958), .A2(g9670), .ZN(g23830) );
AND2_X4 U_g23831 ( .A1(g22962), .A2(g9673), .ZN(g23831) );
AND2_X4 U_g23842 ( .A1(g18207), .A2(g23041), .ZN(g23842) );
AND2_X4 U_g23843 ( .A1(g22966), .A2(g9734), .ZN(g23843) );
AND2_X4 U_g23848 ( .A1(g18226), .A2(g23045), .ZN(g23848) );
AND2_X4 U_g23849 ( .A1(g22771), .A2(g17868), .ZN(g23849) );
AND2_X4 U_g23851 ( .A1(g7329), .A2(g23048), .ZN(g23851) );
AND2_X4 U_g23852 ( .A1(g19179), .A2(g22696), .ZN(g23852) );
AND2_X4 U_g23854 ( .A1(g18265), .A2(g23049), .ZN(g23854) );
AND2_X4 U_g23855 ( .A1(g22954), .A2(g9767), .ZN(g23855) );
AND2_X4 U_g23857 ( .A1(g14263), .A2(g23056), .ZN(g23857) );
AND2_X4 U_g23859 ( .A1(g22958), .A2(g9787), .ZN(g23859) );
AND2_X4 U_g23860 ( .A1(g22962), .A2(g9790), .ZN(g23860) );
AND2_X4 U_g23864 ( .A1(g18297), .A2(g23057), .ZN(g23864) );
AND2_X4 U_g23865 ( .A1(g22966), .A2(g9816), .ZN(g23865) );
AND2_X4 U_g23866 ( .A1(g22971), .A2(g9819), .ZN(g23866) );
AND2_X4 U_g23877 ( .A1(g18314), .A2(g23060), .ZN(g23877) );
AND2_X4 U_g23878 ( .A1(g22975), .A2(g9880), .ZN(g23878) );
AND2_X4 U_g23886 ( .A1(g18341), .A2(g23064), .ZN(g23886) );
AND2_X4 U_g23888 ( .A1(g18358), .A2(g23069), .ZN(g23888) );
AND2_X4 U_g23889 ( .A1(g22962), .A2(g9913), .ZN(g23889) );
AND2_X4 U_g23891 ( .A1(g14385), .A2(g23074), .ZN(g23891) );
AND2_X4 U_g23893 ( .A1(g22966), .A2(g9933), .ZN(g23893) );
AND2_X4 U_g23894 ( .A1(g22971), .A2(g9936), .ZN(g23894) );
AND2_X4 U_g23898 ( .A1(g18390), .A2(g23075), .ZN(g23898) );
AND2_X4 U_g23899 ( .A1(g22975), .A2(g9962), .ZN(g23899) );
AND2_X4 U_g23900 ( .A1(g22980), .A2(g9965), .ZN(g23900) );
AND2_X4 U_g23904 ( .A1(g3010), .A2(g22750), .ZN(g23904) );
AND2_X4 U_g23907 ( .A1(g18436), .A2(g23079), .ZN(g23907) );
AND2_X4 U_g23909 ( .A1(g18453), .A2(g23082), .ZN(g23909) );
AND2_X4 U_g23910 ( .A1(g22971), .A2(g10067), .ZN(g23910) );
AND2_X4 U_g23912 ( .A1(g14497), .A2(g23087), .ZN(g23912) );
AND2_X4 U_g23914 ( .A1(g22975), .A2(g10087), .ZN(g23914) );
AND2_X4 U_g23915 ( .A1(g22980), .A2(g10090), .ZN(g23915) );
AND2_X4 U_g23917 ( .A1(g7545), .A2(g23088), .ZN(g23917) );
AND2_X4 U_g23939 ( .A1(g18509), .A2(g23095), .ZN(g23939) );
AND2_X4 U_g23941 ( .A1(g18526), .A2(g23098), .ZN(g23941) );
AND2_X4 U_g23942 ( .A1(g22980), .A2(g10176), .ZN(g23942) );
AND2_X4 U_g23944 ( .A1(g7570), .A2(g23103), .ZN(g23944) );
AND2_X4 U_g23971 ( .A1(g18573), .A2(g23112), .ZN(g23971) );
AND2_X4 U_g23972 ( .A1(g2903), .A2(g23115), .ZN(g23972) );
AND2_X4 U_g24029 ( .A1(g2900), .A2(g22903), .ZN(g24029) );
AND2_X4 U_g24211 ( .A1(g22014), .A2(g10969), .ZN(g24211) );
AND2_X4 U_g24217 ( .A1(g22825), .A2(g10999), .ZN(g24217) );
AND2_X4 U_g24221 ( .A1(g22979), .A2(g11042), .ZN(g24221) );
AND2_X4 U_g24224 ( .A1(g22219), .A2(g11045), .ZN(g24224) );
AND2_X4 U_g24229 ( .A1(g22232), .A2(g11105), .ZN(g24229) );
AND2_X4 U_g24236 ( .A1(g22243), .A2(g11157), .ZN(g24236) );
AND2_X4 U_g24241 ( .A1(g22259), .A2(g11228), .ZN(g24241) );
AND2_X4 U_g24246 ( .A1(g21982), .A2(g11291), .ZN(g24246) );
AND2_X4 U_g24247 ( .A1(g22551), .A2(g11297), .ZN(g24247) );
AND2_X4 U_g24253 ( .A1(g21995), .A2(g11370), .ZN(g24253) );
AND2_X4 U_g24256 ( .A1(g22003), .A2(g11438), .ZN(g24256) );
AND3_X4 U_g24427 ( .A1(g17086), .A2(g24134), .A3(g13626), .ZN(g24427) );
AND2_X4 U_g24429 ( .A1(g24115), .A2(g13614), .ZN(g24429) );
AND3_X4 U_g24431 ( .A1(g17124), .A2(g24153), .A3(g13637), .ZN(g24431) );
AND3_X4 U_g24432 ( .A1(g14642), .A2(g15904), .A3(g24115), .ZN(g24432) );
AND2_X4 U_g24433 ( .A1(g24134), .A2(g13626), .ZN(g24433) );
AND3_X4 U_g24435 ( .A1(g17151), .A2(g24168), .A3(g13649), .ZN(g24435) );
AND3_X4 U_g24436 ( .A1(g14669), .A2(g15933), .A3(g24134), .ZN(g24436) );
AND2_X4 U_g24437 ( .A1(g24153), .A2(g13637), .ZN(g24437) );
AND3_X4 U_g24439 ( .A1(g14703), .A2(g15962), .A3(g24153), .ZN(g24439) );
AND2_X4 U_g24440 ( .A1(g24168), .A2(g13649), .ZN(g24440) );
AND3_X4 U_g24441 ( .A1(g14737), .A2(g15981), .A3(g24168), .ZN(g24441) );
AND3_X4 U_g24478 ( .A1(g23545), .A2(g21119), .A3(g21227), .ZN(g24478) );
AND3_X4 U_g24529 ( .A1(g19933), .A2(g17896), .A3(g23403), .ZN(g24529) );
AND3_X4 U_g24540 ( .A1(g18548), .A2(g23089), .A3(g23403), .ZN(g24540) );
AND3_X4 U_g24541 ( .A1(g23420), .A2(g17896), .A3(g23052), .ZN(g24541) );
AND3_X4 U_g24542 ( .A1(g19950), .A2(g18007), .A3(g23410), .ZN(g24542) );
AND3_X4 U_g24550 ( .A1(g18548), .A2(g23420), .A3(g19948), .ZN(g24550) );
AND3_X4 U_g24552 ( .A1(g18598), .A2(g23107), .A3(g23410), .ZN(g24552) );
AND3_X4 U_g24553 ( .A1(g23429), .A2(g18007), .A3(g23071), .ZN(g24553) );
AND3_X4 U_g24554 ( .A1(g19977), .A2(g18124), .A3(g23415), .ZN(g24554) );
AND2_X4 U_g24559 ( .A1(g79), .A2(g23448), .ZN(g24559) );
AND3_X4 U_g24561 ( .A1(g18598), .A2(g23429), .A3(g19975), .ZN(g24561) );
AND3_X4 U_g24563 ( .A1(g18630), .A2(g23120), .A3(g23415), .ZN(g24563) );
AND3_X4 U_g24564 ( .A1(g23435), .A2(g18124), .A3(g23084), .ZN(g24564) );
AND3_X4 U_g24565 ( .A1(g20007), .A2(g18240), .A3(g23424), .ZN(g24565) );
AND2_X4 U_g24569 ( .A1(g767), .A2(g23455), .ZN(g24569) );
AND3_X4 U_g24571 ( .A1(g18630), .A2(g23435), .A3(g20005), .ZN(g24571) );
AND3_X4 U_g24573 ( .A1(g18639), .A2(g23129), .A3(g23424), .ZN(g24573) );
AND3_X4 U_g24574 ( .A1(g23441), .A2(g18240), .A3(g23100), .ZN(g24574) );
AND2_X4 U_g24578 ( .A1(g1453), .A2(g23464), .ZN(g24578) );
AND3_X4 U_g24580 ( .A1(g18639), .A2(g23441), .A3(g20043), .ZN(g24580) );
AND2_X4 U_g24585 ( .A1(g2147), .A2(g23473), .ZN(g24585) );
AND2_X4 U_g24590 ( .A1(g23486), .A2(g23478), .ZN(g24590) );
AND2_X4 U_g24591 ( .A1(g83), .A2(g23853), .ZN(g24591) );
AND2_X4 U_g24595 ( .A1(g23502), .A2(g23489), .ZN(g24595) );
AND2_X4 U_g24596 ( .A1(g771), .A2(g23887), .ZN(g24596) );
AND2_X4 U_g24603 ( .A1(g23518), .A2(g23505), .ZN(g24603) );
AND2_X4 U_g24604 ( .A1(g1457), .A2(g23908), .ZN(g24604) );
AND2_X4 U_g24610 ( .A1(g23533), .A2(g23521), .ZN(g24610) );
AND2_X4 U_g24611 ( .A1(g2151), .A2(g23940), .ZN(g24611) );
AND2_X4 U_g24644 ( .A1(g17203), .A2(g24115), .ZN(g24644) );
AND2_X4 U_g24664 ( .A1(g17208), .A2(g24134), .ZN(g24664) );
AND2_X4 U_g24676 ( .A1(g13568), .A2(g24115), .ZN(g24676) );
AND2_X4 U_g24683 ( .A1(g17214), .A2(g24153), .ZN(g24683) );
AND2_X4 U_g24695 ( .A1(g13576), .A2(g24134), .ZN(g24695) );
AND2_X4 U_g24700 ( .A1(g17217), .A2(g24168), .ZN(g24700) );
AND2_X4 U_g24712 ( .A1(g13585), .A2(g24153), .ZN(g24712) );
AND2_X4 U_g24723 ( .A1(g13605), .A2(g24168), .ZN(g24723) );
AND2_X4 U_g24745 ( .A1(g15454), .A2(g24096), .ZN(g24745) );
AND2_X4 U_g24746 ( .A1(g15454), .A2(g24098), .ZN(g24746) );
AND2_X4 U_g24747 ( .A1(g9427), .A2(g24099), .ZN(g24747) );
AND2_X4 U_g24748 ( .A1(g672), .A2(g24101), .ZN(g24748) );
AND2_X4 U_g24749 ( .A1(g15540), .A2(g24102), .ZN(g24749) );
AND2_X4 U_g24750 ( .A1(g15454), .A2(g24104), .ZN(g24750) );
AND2_X4 U_g24751 ( .A1(g9427), .A2(g24105), .ZN(g24751) );
AND2_X4 U_g24752 ( .A1(g9507), .A2(g24106), .ZN(g24752) );
AND2_X4 U_g24754 ( .A1(g15540), .A2(g24107), .ZN(g24754) );
AND2_X4 U_g24755 ( .A1(g9569), .A2(g24108), .ZN(g24755) );
AND2_X4 U_g24757 ( .A1(g1358), .A2(g24110), .ZN(g24757) );
AND2_X4 U_g24758 ( .A1(g15618), .A2(g24111), .ZN(g24758) );
AND2_X4 U_g24759 ( .A1(g21825), .A2(g23885), .ZN(g24759) );
AND2_X4 U_g24760 ( .A1(g9427), .A2(g24112), .ZN(g24760) );
AND2_X4 U_g24761 ( .A1(g9507), .A2(g24113), .ZN(g24761) );
AND2_X4 U_g24762 ( .A1(g12876), .A2(g24114), .ZN(g24762) );
AND2_X4 U_g24767 ( .A1(g15540), .A2(g24121), .ZN(g24767) );
AND2_X4 U_g24768 ( .A1(g9569), .A2(g24122), .ZN(g24768) );
AND2_X4 U_g24769 ( .A1(g9649), .A2(g24123), .ZN(g24769) );
AND2_X4 U_g24772 ( .A1(g15618), .A2(g24124), .ZN(g24772) );
AND2_X4 U_g24773 ( .A1(g9711), .A2(g24125), .ZN(g24773) );
AND2_X4 U_g24774 ( .A1(g2052), .A2(g24127), .ZN(g24774) );
AND2_X4 U_g24775 ( .A1(g15694), .A2(g24128), .ZN(g24775) );
AND2_X4 U_g24776 ( .A1(g9507), .A2(g24129), .ZN(g24776) );
AND2_X4 U_g24777 ( .A1(g12876), .A2(g24130), .ZN(g24777) );
AND2_X4 U_g24779 ( .A1(g9569), .A2(g24131), .ZN(g24779) );
AND2_X4 U_g24780 ( .A1(g9649), .A2(g24132), .ZN(g24780) );
AND2_X4 U_g24781 ( .A1(g12916), .A2(g24133), .ZN(g24781) );
AND2_X4 U_g24788 ( .A1(g15618), .A2(g24140), .ZN(g24788) );
AND2_X4 U_g24789 ( .A1(g9711), .A2(g24141), .ZN(g24789) );
AND2_X4 U_g24790 ( .A1(g9795), .A2(g24142), .ZN(g24790) );
AND2_X4 U_g24792 ( .A1(g15694), .A2(g24143), .ZN(g24792) );
AND2_X4 U_g24793 ( .A1(g9857), .A2(g24144), .ZN(g24793) );
AND2_X4 U_g24794 ( .A1(g2746), .A2(g24146), .ZN(g24794) );
AND2_X4 U_g24795 ( .A1(g12017), .A2(g24232), .ZN(g24795) );
AND2_X4 U_g24796 ( .A1(g12876), .A2(g24147), .ZN(g24796) );
AND2_X4 U_g24798 ( .A1(g9649), .A2(g24148), .ZN(g24798) );
AND2_X4 U_g24799 ( .A1(g12916), .A2(g24149), .ZN(g24799) );
AND2_X4 U_g24802 ( .A1(g9711), .A2(g24150), .ZN(g24802) );
AND2_X4 U_g24803 ( .A1(g9795), .A2(g24151), .ZN(g24803) );
AND2_X4 U_g24804 ( .A1(g12945), .A2(g24152), .ZN(g24804) );
AND2_X4 U_g24809 ( .A1(g15694), .A2(g24159), .ZN(g24809) );
AND2_X4 U_g24810 ( .A1(g9857), .A2(g24160), .ZN(g24810) );
AND2_X4 U_g24811 ( .A1(g9941), .A2(g24161), .ZN(g24811) );
AND2_X4 U_g24813 ( .A1(g21825), .A2(g23905), .ZN(g24813) );
AND2_X4 U_g24818 ( .A1(g12916), .A2(g24162), .ZN(g24818) );
AND2_X4 U_g24821 ( .A1(g9795), .A2(g24163), .ZN(g24821) );
AND2_X4 U_g24822 ( .A1(g12945), .A2(g24164), .ZN(g24822) );
AND2_X4 U_g24824 ( .A1(g9857), .A2(g24165), .ZN(g24824) );
AND2_X4 U_g24825 ( .A1(g9941), .A2(g24166), .ZN(g24825) );
AND2_X4 U_g24826 ( .A1(g12974), .A2(g24167), .ZN(g24826) );
AND2_X4 U_g24831 ( .A1(g24100), .A2(g20401), .ZN(g24831) );
AND2_X4 U_g24838 ( .A1(g12945), .A2(g24175), .ZN(g24838) );
AND2_X4 U_g24840 ( .A1(g9941), .A2(g24176), .ZN(g24840) );
AND2_X4 U_g24841 ( .A1(g12974), .A2(g24177), .ZN(g24841) );
AND2_X4 U_g24843 ( .A1(g21825), .A2(g23918), .ZN(g24843) );
AND2_X4 U_g24846 ( .A1(g24109), .A2(g20426), .ZN(g24846) );
AND2_X4 U_g24853 ( .A1(g12974), .A2(g24180), .ZN(g24853) );
AND2_X4 U_g24855 ( .A1(g18174), .A2(g23731), .ZN(g24855) );
AND2_X4 U_g24858 ( .A1(g24047), .A2(g18873), .ZN(g24858) );
AND2_X4 U_g24861 ( .A1(g24126), .A2(g20448), .ZN(g24861) );
AND2_X4 U_g24867 ( .A1(g666), .A2(g23779), .ZN(g24867) );
AND2_X4 U_g24869 ( .A1(g24047), .A2(g18894), .ZN(g24869) );
AND2_X4 U_g24870 ( .A1(g18281), .A2(g23786), .ZN(g24870) );
AND2_X4 U_g24874 ( .A1(g24060), .A2(g18899), .ZN(g24874) );
AND2_X4 U_g24876 ( .A1(g24145), .A2(g20467), .ZN(g24876) );
AND2_X4 U_g24878 ( .A1(g19830), .A2(g24210), .ZN(g24878) );
AND2_X4 U_g24881 ( .A1(g24047), .A2(g18912), .ZN(g24881) );
AND2_X4 U_g24882 ( .A1(g1352), .A2(g23832), .ZN(g24882) );
AND2_X4 U_g24884 ( .A1(g24060), .A2(g18917), .ZN(g24884) );
AND2_X4 U_g24885 ( .A1(g18374), .A2(g23839), .ZN(g24885) );
AND2_X4 U_g24888 ( .A1(g24073), .A2(g18922), .ZN(g24888) );
AND2_X4 U_g24898 ( .A1(g24060), .A2(g18931), .ZN(g24898) );
AND2_X4 U_g24899 ( .A1(g2046), .A2(g23867), .ZN(g24899) );
AND2_X4 U_g24901 ( .A1(g24073), .A2(g18936), .ZN(g24901) );
AND2_X4 U_g24902 ( .A1(g18469), .A2(g23874), .ZN(g24902) );
AND2_X4 U_g24905 ( .A1(g24084), .A2(g18941), .ZN(g24905) );
AND2_X4 U_g24906 ( .A1(g18886), .A2(g23879), .ZN(g24906) );
AND2_X4 U_g24907 ( .A1(g7466), .A2(g24220), .ZN(g24907) );
AND2_X4 U_g24908 ( .A1(g7342), .A2(g23882), .ZN(g24908) );
AND2_X4 U_g24921 ( .A1(g24073), .A2(g18951), .ZN(g24921) );
AND2_X4 U_g24922 ( .A1(g2740), .A2(g23901), .ZN(g24922) );
AND2_X4 U_g24924 ( .A1(g24084), .A2(g18956), .ZN(g24924) );
AND2_X4 U_g24938 ( .A1(g24084), .A2(g18967), .ZN(g24938) );
AND2_X4 U_g24964 ( .A1(g7595), .A2(g24251), .ZN(g24964) );
AND2_X4 U_g24974 ( .A1(g7600), .A2(g24030), .ZN(g24974) );
AND2_X4 U_g25086 ( .A1(g23444), .A2(g10880), .ZN(g25086) );
AND2_X4 U_g25102 ( .A1(g23444), .A2(g10915), .ZN(g25102) );
AND2_X4 U_g25117 ( .A1(g23444), .A2(g10974), .ZN(g25117) );
AND3_X4 U_g25128 ( .A1(g17051), .A2(g24115), .A3(g13614), .ZN(g25128) );
AND2_X4 U_g25178 ( .A1(g24623), .A2(g20634), .ZN(g25178) );
AND2_X4 U_g25181 ( .A1(g24636), .A2(g20673), .ZN(g25181) );
AND2_X4 U_g25182 ( .A1(g24681), .A2(g20676), .ZN(g25182) );
AND2_X4 U_g25184 ( .A1(g24694), .A2(g20735), .ZN(g25184) );
AND2_X4 U_g25187 ( .A1(g24633), .A2(g16608), .ZN(g25187) );
AND2_X4 U_g25188 ( .A1(g24652), .A2(g20763), .ZN(g25188) );
AND2_X4 U_g25192 ( .A1(g24711), .A2(g20790), .ZN(g25192) );
AND2_X4 U_g25193 ( .A1(g24653), .A2(g16626), .ZN(g25193) );
AND2_X4 U_g25196 ( .A1(g24672), .A2(g16640), .ZN(g25196) );
AND2_X4 U_g25198 ( .A1(g24691), .A2(g16651), .ZN(g25198) );
AND2_X4 U_g25269 ( .A1(g24648), .A2(g8700), .ZN(g25269) );
AND2_X4 U_g25277 ( .A1(g24648), .A2(g8714), .ZN(g25277) );
AND2_X4 U_g25278 ( .A1(g24668), .A2(g8719), .ZN(g25278) );
AND2_X4 U_g25281 ( .A1(g5606), .A2(g24815), .ZN(g25281) );
AND2_X4 U_g25282 ( .A1(g24648), .A2(g8748), .ZN(g25282) );
AND2_X4 U_g25286 ( .A1(g24668), .A2(g8752), .ZN(g25286) );
AND2_X4 U_g25287 ( .A1(g24687), .A2(g8757), .ZN(g25287) );
AND2_X4 U_g25289 ( .A1(g5631), .A2(g24834), .ZN(g25289) );
AND2_X4 U_g25290 ( .A1(g24668), .A2(g8771), .ZN(g25290) );
AND2_X4 U_g25294 ( .A1(g24687), .A2(g8775), .ZN(g25294) );
AND2_X4 U_g25295 ( .A1(g24704), .A2(g8780), .ZN(g25295) );
AND2_X4 U_g25299 ( .A1(g5659), .A2(g24850), .ZN(g25299) );
AND2_X4 U_g25300 ( .A1(g24687), .A2(g8794), .ZN(g25300) );
AND2_X4 U_g25304 ( .A1(g24704), .A2(g8798), .ZN(g25304) );
AND2_X4 U_g25309 ( .A1(g5697), .A2(g24864), .ZN(g25309) );
AND2_X4 U_g25310 ( .A1(g24704), .A2(g8813), .ZN(g25310) );
AND3_X4 U_g25318 ( .A1(g24682), .A2(g19358), .A3(g19335), .ZN(g25318) );
AND2_X4 U_g25321 ( .A1(g25075), .A2(g9669), .ZN(g25321) );
AND2_X4 U_g25328 ( .A1(g24644), .A2(g17892), .ZN(g25328) );
AND2_X4 U_g25334 ( .A1(g24644), .A2(g17984), .ZN(g25334) );
AND2_X4 U_g25337 ( .A1(g24664), .A2(g18003), .ZN(g25337) );
AND2_X4 U_g25342 ( .A1(g5851), .A2(g24600), .ZN(g25342) );
AND2_X4 U_g25346 ( .A1(g24644), .A2(g18084), .ZN(g25346) );
AND2_X4 U_g25348 ( .A1(g24664), .A2(g18101), .ZN(g25348) );
AND2_X4 U_g25351 ( .A1(g24683), .A2(g18120), .ZN(g25351) );
AND2_X4 U_g25356 ( .A1(g5898), .A2(g24607), .ZN(g25356) );
AND2_X4 U_g25360 ( .A1(g24664), .A2(g18200), .ZN(g25360) );
AND2_X4 U_g25362 ( .A1(g24683), .A2(g18217), .ZN(g25362) );
AND2_X4 U_g25365 ( .A1(g24700), .A2(g18236), .ZN(g25365) );
AND2_X4 U_g25371 ( .A1(g5937), .A2(g24619), .ZN(g25371) );
AND2_X4 U_g25375 ( .A1(g24683), .A2(g18307), .ZN(g25375) );
AND2_X4 U_g25377 ( .A1(g24700), .A2(g18324), .ZN(g25377) );
AND2_X4 U_g25388 ( .A1(g5971), .A2(g24630), .ZN(g25388) );
AND2_X4 U_g25392 ( .A1(g24700), .A2(g18400), .ZN(g25392) );
AND2_X4 U_g25453 ( .A1(g6142), .A2(g24763), .ZN(g25453) );
AND2_X4 U_g25457 ( .A1(g6163), .A2(g24784), .ZN(g25457) );
AND2_X4 U_g25461 ( .A1(g6190), .A2(g24805), .ZN(g25461) );
AND2_X4 U_g25466 ( .A1(g6222), .A2(g24827), .ZN(g25466) );
AND2_X4 U_g25470 ( .A1(g24479), .A2(g20400), .ZN(g25470) );
AND2_X4 U_g25475 ( .A1(g14148), .A2(g25087), .ZN(g25475) );
AND2_X4 U_g25482 ( .A1(g24480), .A2(g17567), .ZN(g25482) );
AND2_X4 U_g25483 ( .A1(g24481), .A2(g20421), .ZN(g25483) );
AND2_X4 U_g25487 ( .A1(g24485), .A2(g20425), .ZN(g25487) );
AND2_X4 U_g25505 ( .A1(g6707), .A2(g25094), .ZN(g25505) );
AND2_X4 U_g25506 ( .A1(g14263), .A2(g25095), .ZN(g25506) );
AND2_X4 U_g25513 ( .A1(g24487), .A2(g17664), .ZN(g25513) );
AND2_X4 U_g25514 ( .A1(g24488), .A2(g20443), .ZN(g25514) );
AND2_X4 U_g25518 ( .A1(g24489), .A2(g20447), .ZN(g25518) );
AND2_X4 U_g25552 ( .A1(g7009), .A2(g25104), .ZN(g25552) );
AND2_X4 U_g25553 ( .A1(g14385), .A2(g25105), .ZN(g25553) );
AND2_X4 U_g25560 ( .A1(g24494), .A2(g17764), .ZN(g25560) );
AND2_X4 U_g25561 ( .A1(g24495), .A2(g20462), .ZN(g25561) );
AND2_X4 U_g25565 ( .A1(g24496), .A2(g20466), .ZN(g25565) );
AND2_X4 U_g25618 ( .A1(g7259), .A2(g25110), .ZN(g25618) );
AND2_X4 U_g25619 ( .A1(g14497), .A2(g25111), .ZN(g25619) );
AND2_X4 U_g25626 ( .A1(g24504), .A2(g17865), .ZN(g25626) );
AND2_X4 U_g25627 ( .A1(g24505), .A2(g20477), .ZN(g25627) );
AND2_X4 U_g25628 ( .A1(g21008), .A2(g25115), .ZN(g25628) );
AND2_X4 U_g25629 ( .A1(g3024), .A2(g25116), .ZN(g25629) );
AND2_X4 U_g25697 ( .A1(g7455), .A2(g25120), .ZN(g25697) );
AND2_X4 U_g25881 ( .A1(g2908), .A2(g25126), .ZN(g25881) );
AND2_X4 U_g25951 ( .A1(g24800), .A2(g13670), .ZN(g25951) );
AND2_X4 U_g25953 ( .A1(g24783), .A2(g13699), .ZN(g25953) );
AND2_X4 U_g25957 ( .A1(g24782), .A2(g11869), .ZN(g25957) );
AND2_X4 U_g25961 ( .A1(g24770), .A2(g11901), .ZN(g25961) );
AND2_X4 U_g25963 ( .A1(g24756), .A2(g11944), .ZN(g25963) );
AND2_X4 U_g25968 ( .A1(g24871), .A2(g11986), .ZN(g25968) );
AND2_X4 U_g25972 ( .A1(g24859), .A2(g12042), .ZN(g25972) );
AND2_X4 U_g25973 ( .A1(g24847), .A2(g13838), .ZN(g25973) );
AND2_X4 U_g25975 ( .A1(g24606), .A2(g21917), .ZN(g25975) );
AND2_X4 U_g25977 ( .A1(g24845), .A2(g12089), .ZN(g25977) );
AND2_X4 U_g25978 ( .A1(g24836), .A2(g13850), .ZN(g25978) );
AND2_X4 U_g25980 ( .A1(g24663), .A2(g21928), .ZN(g25980) );
AND2_X4 U_g25981 ( .A1(g24819), .A2(g13858), .ZN(g25981) );
AND2_X4 U_g26023 ( .A1(g25422), .A2(g24912), .ZN(g26023) );
AND2_X4 U_g26024 ( .A1(g25301), .A2(g21102), .ZN(g26024) );
AND2_X4 U_g26026 ( .A1(g25431), .A2(g24929), .ZN(g26026) );
AND2_X4 U_g26027 ( .A1(g25418), .A2(g22271), .ZN(g26027) );
AND2_X4 U_g26028 ( .A1(g25438), .A2(g24941), .ZN(g26028) );
AND2_X4 U_g26029 ( .A1(g25445), .A2(g24952), .ZN(g26029) );
AND2_X4 U_g26030 ( .A1(g25429), .A2(g22304), .ZN(g26030) );
AND2_X4 U_g26032 ( .A1(g25379), .A2(g19415), .ZN(g26032) );
AND2_X4 U_g26033 ( .A1(g25395), .A2(g19452), .ZN(g26033) );
AND2_X4 U_g26034 ( .A1(g25405), .A2(g19479), .ZN(g26034) );
AND2_X4 U_g26035 ( .A1(g25523), .A2(g19483), .ZN(g26035) );
AND2_X4 U_g26036 ( .A1(g25413), .A2(g19502), .ZN(g26036) );
AND2_X4 U_g26038 ( .A1(g25589), .A2(g19504), .ZN(g26038) );
AND2_X4 U_g26039 ( .A1(g25668), .A2(g19523), .ZN(g26039) );
AND2_X4 U_g26040 ( .A1(g25745), .A2(g19533), .ZN(g26040) );
AND2_X4 U_g26051 ( .A1(g70), .A2(g25296), .ZN(g26051) );
AND2_X4 U_g26052 ( .A1(g25941), .A2(g21087), .ZN(g26052) );
AND2_X4 U_g26053 ( .A1(g758), .A2(g25306), .ZN(g26053) );
AND2_X4 U_g26054 ( .A1(g25944), .A2(g21099), .ZN(g26054) );
AND2_X4 U_g26060 ( .A1(g25943), .A2(g21108), .ZN(g26060) );
AND2_X4 U_g26061 ( .A1(g1444), .A2(g25315), .ZN(g26061) );
AND2_X4 U_g26062 ( .A1(g25947), .A2(g21113), .ZN(g26062) );
AND2_X4 U_g26067 ( .A1(g25946), .A2(g21125), .ZN(g26067) );
AND2_X4 U_g26068 ( .A1(g2138), .A2(g25324), .ZN(g26068) );
AND2_X4 U_g26069 ( .A1(g25949), .A2(g21130), .ZN(g26069) );
AND2_X4 U_g26074 ( .A1(g25948), .A2(g21144), .ZN(g26074) );
AND2_X4 U_g26075 ( .A1(g74), .A2(g25698), .ZN(g26075) );
AND2_X4 U_g26080 ( .A1(g25950), .A2(g21164), .ZN(g26080) );
AND2_X4 U_g26082 ( .A1(g762), .A2(g25771), .ZN(g26082) );
AND2_X4 U_g26085 ( .A1(g1448), .A2(g25825), .ZN(g26085) );
AND2_X4 U_g26091 ( .A1(g2142), .A2(g25860), .ZN(g26091) );
AND2_X4 U_g26157 ( .A1(g21825), .A2(g25630), .ZN(g26157) );
AND2_X4 U_g26158 ( .A1(g679), .A2(g25937), .ZN(g26158) );
AND2_X4 U_g26163 ( .A1(g1365), .A2(g25939), .ZN(g26163) );
AND2_X4 U_g26166 ( .A1(g686), .A2(g25454), .ZN(g26166) );
AND2_X4 U_g26171 ( .A1(g2059), .A2(g25942), .ZN(g26171) );
AND2_X4 U_g26186 ( .A1(g1372), .A2(g25458), .ZN(g26186) );
AND2_X4 U_g26188 ( .A1(g2753), .A2(g25945), .ZN(g26188) );
AND2_X4 U_g26207 ( .A1(g2066), .A2(g25463), .ZN(g26207) );
AND2_X4 U_g26212 ( .A1(g4217), .A2(g25467), .ZN(g26212) );
AND2_X4 U_g26213 ( .A1(g25895), .A2(g9306), .ZN(g26213) );
AND2_X4 U_g26231 ( .A1(g2760), .A2(g25472), .ZN(g26231) );
AND2_X4 U_g26233 ( .A1(g4340), .A2(g25476), .ZN(g26233) );
AND2_X4 U_g26234 ( .A1(g4343), .A2(g25479), .ZN(g26234) );
AND2_X4 U_g26235 ( .A1(g25895), .A2(g9368), .ZN(g26235) );
AND2_X4 U_g26236 ( .A1(g25899), .A2(g9371), .ZN(g26236) );
AND2_X4 U_g26243 ( .A1(g4372), .A2(g25484), .ZN(g26243) );
AND2_X4 U_g26244 ( .A1(g25903), .A2(g9387), .ZN(g26244) );
AND2_X4 U_g26257 ( .A1(g4465), .A2(g25493), .ZN(g26257) );
AND2_X4 U_g26258 ( .A1(g4468), .A2(g25496), .ZN(g26258) );
AND2_X4 U_g26259 ( .A1(g4471), .A2(g25499), .ZN(g26259) );
AND2_X4 U_g26260 ( .A1(g25254), .A2(g17649), .ZN(g26260) );
AND2_X4 U_g26261 ( .A1(g25895), .A2(g9443), .ZN(g26261) );
AND2_X4 U_g26262 ( .A1(g25899), .A2(g9446), .ZN(g26262) );
AND2_X4 U_g26263 ( .A1(g4476), .A2(g25502), .ZN(g26263) );
AND2_X4 U_g26268 ( .A1(g4509), .A2(g25507), .ZN(g26268) );
AND2_X4 U_g26269 ( .A1(g4512), .A2(g25510), .ZN(g26269) );
AND2_X4 U_g26270 ( .A1(g25903), .A2(g9465), .ZN(g26270) );
AND2_X4 U_g26271 ( .A1(g25907), .A2(g9468), .ZN(g26271) );
AND2_X4 U_g26278 ( .A1(g4541), .A2(g25515), .ZN(g26278) );
AND2_X4 U_g26279 ( .A1(g25911), .A2(g9484), .ZN(g26279) );
AND2_X4 U_g26288 ( .A1(g4592), .A2(g25524), .ZN(g26288) );
AND2_X4 U_g26289 ( .A1(g4595), .A2(g25527), .ZN(g26289) );
AND2_X4 U_g26290 ( .A1(g4598), .A2(g25530), .ZN(g26290) );
AND2_X4 U_g26291 ( .A1(g25899), .A2(g9524), .ZN(g26291) );
AND2_X4 U_g26292 ( .A1(g4603), .A2(g25533), .ZN(g26292) );
AND2_X4 U_g26293 ( .A1(g4606), .A2(g25536), .ZN(g26293) );
AND2_X4 U_g26298 ( .A1(g4641), .A2(g25540), .ZN(g26298) );
AND2_X4 U_g26299 ( .A1(g4644), .A2(g25543), .ZN(g26299) );
AND2_X4 U_g26300 ( .A1(g4647), .A2(g25546), .ZN(g26300) );
AND2_X4 U_g26301 ( .A1(g25258), .A2(g17749), .ZN(g26301) );
AND2_X4 U_g26302 ( .A1(g25903), .A2(g9585), .ZN(g26302) );
AND2_X4 U_g26303 ( .A1(g25907), .A2(g9588), .ZN(g26303) );
AND2_X4 U_g26307 ( .A1(g4652), .A2(g25549), .ZN(g26307) );
AND2_X4 U_g26309 ( .A1(g4685), .A2(g25554), .ZN(g26309) );
AND2_X4 U_g26310 ( .A1(g4688), .A2(g25557), .ZN(g26310) );
AND2_X4 U_g26311 ( .A1(g25911), .A2(g9607), .ZN(g26311) );
AND2_X4 U_g26312 ( .A1(g25915), .A2(g9610), .ZN(g26312) );
AND2_X4 U_g26316 ( .A1(g4717), .A2(g25562), .ZN(g26316) );
AND2_X4 U_g26317 ( .A1(g25919), .A2(g9626), .ZN(g26317) );
AND2_X4 U_g26318 ( .A1(g4737), .A2(g25573), .ZN(g26318) );
AND2_X4 U_g26319 ( .A1(g4740), .A2(g25576), .ZN(g26319) );
AND2_X4 U_g26324 ( .A1(g4743), .A2(g25579), .ZN(g26324) );
AND2_X4 U_g26325 ( .A1(g4746), .A2(g25582), .ZN(g26325) );
AND2_X4 U_g26326 ( .A1(g4749), .A2(g25585), .ZN(g26326) );
AND2_X4 U_g26332 ( .A1(g4769), .A2(g25590), .ZN(g26332) );
AND2_X4 U_g26333 ( .A1(g4772), .A2(g25593), .ZN(g26333) );
AND2_X4 U_g26334 ( .A1(g4775), .A2(g25596), .ZN(g26334) );
AND2_X4 U_g26335 ( .A1(g25907), .A2(g9666), .ZN(g26335) );
AND2_X4 U_g26339 ( .A1(g4780), .A2(g25599), .ZN(g26339) );
AND2_X4 U_g26340 ( .A1(g4783), .A2(g25602), .ZN(g26340) );
AND2_X4 U_g26342 ( .A1(g4818), .A2(g25606), .ZN(g26342) );
AND2_X4 U_g26343 ( .A1(g4821), .A2(g25609), .ZN(g26343) );
AND2_X4 U_g26344 ( .A1(g4824), .A2(g25612), .ZN(g26344) );
AND2_X4 U_g26345 ( .A1(g25261), .A2(g17850), .ZN(g26345) );
AND2_X4 U_g26346 ( .A1(g25911), .A2(g9727), .ZN(g26346) );
AND2_X4 U_g26347 ( .A1(g25915), .A2(g9730), .ZN(g26347) );
AND2_X4 U_g26348 ( .A1(g4829), .A2(g25615), .ZN(g26348) );
AND2_X4 U_g26350 ( .A1(g4862), .A2(g25620), .ZN(g26350) );
AND2_X4 U_g26351 ( .A1(g4865), .A2(g25623), .ZN(g26351) );
AND2_X4 U_g26352 ( .A1(g25919), .A2(g9749), .ZN(g26352) );
AND2_X4 U_g26353 ( .A1(g25923), .A2(g9752), .ZN(g26353) );
AND2_X4 U_g26357 ( .A1(g4882), .A2(g25634), .ZN(g26357) );
AND2_X4 U_g26361 ( .A1(g4888), .A2(g25637), .ZN(g26361) );
AND2_X4 U_g26362 ( .A1(g4891), .A2(g25640), .ZN(g26362) );
AND2_X4 U_g26363 ( .A1(g4894), .A2(g25643), .ZN(g26363) );
AND2_X4 U_g26365 ( .A1(g4913), .A2(g25652), .ZN(g26365) );
AND2_X4 U_g26366 ( .A1(g4916), .A2(g25655), .ZN(g26366) );
AND2_X4 U_g26371 ( .A1(g4919), .A2(g25658), .ZN(g26371) );
AND2_X4 U_g26372 ( .A1(g4922), .A2(g25661), .ZN(g26372) );
AND2_X4 U_g26373 ( .A1(g4925), .A2(g25664), .ZN(g26373) );
AND2_X4 U_g26379 ( .A1(g4945), .A2(g25669), .ZN(g26379) );
AND2_X4 U_g26380 ( .A1(g4948), .A2(g25672), .ZN(g26380) );
AND2_X4 U_g26381 ( .A1(g4951), .A2(g25675), .ZN(g26381) );
AND2_X4 U_g26382 ( .A1(g25915), .A2(g9812), .ZN(g26382) );
AND2_X4 U_g26383 ( .A1(g4956), .A2(g25678), .ZN(g26383) );
AND2_X4 U_g26384 ( .A1(g4959), .A2(g25681), .ZN(g26384) );
AND2_X4 U_g26386 ( .A1(g4994), .A2(g25685), .ZN(g26386) );
AND2_X4 U_g26387 ( .A1(g4997), .A2(g25688), .ZN(g26387) );
AND2_X4 U_g26388 ( .A1(g5000), .A2(g25691), .ZN(g26388) );
AND2_X4 U_g26389 ( .A1(g25264), .A2(g17962), .ZN(g26389) );
AND2_X4 U_g26390 ( .A1(g25919), .A2(g9873), .ZN(g26390) );
AND2_X4 U_g26391 ( .A1(g25923), .A2(g9876), .ZN(g26391) );
AND2_X4 U_g26392 ( .A1(g5005), .A2(g25694), .ZN(g26392) );
AND2_X4 U_g26396 ( .A1(g5027), .A2(g25700), .ZN(g26396) );
AND2_X4 U_g26397 ( .A1(g5030), .A2(g25703), .ZN(g26397) );
AND2_X4 U_g26400 ( .A1(g5041), .A2(g25711), .ZN(g26400) );
AND2_X4 U_g26404 ( .A1(g5047), .A2(g25714), .ZN(g26404) );
AND2_X4 U_g26405 ( .A1(g5050), .A2(g25717), .ZN(g26405) );
AND2_X4 U_g26406 ( .A1(g5053), .A2(g25720), .ZN(g26406) );
AND2_X4 U_g26408 ( .A1(g5072), .A2(g25729), .ZN(g26408) );
AND2_X4 U_g26409 ( .A1(g5075), .A2(g25732), .ZN(g26409) );
AND2_X4 U_g26414 ( .A1(g5078), .A2(g25735), .ZN(g26414) );
AND2_X4 U_g26415 ( .A1(g5081), .A2(g25738), .ZN(g26415) );
AND2_X4 U_g26416 ( .A1(g5084), .A2(g25741), .ZN(g26416) );
AND2_X4 U_g26422 ( .A1(g5104), .A2(g25746), .ZN(g26422) );
AND2_X4 U_g26423 ( .A1(g5107), .A2(g25749), .ZN(g26423) );
AND2_X4 U_g26424 ( .A1(g5110), .A2(g25752), .ZN(g26424) );
AND2_X4 U_g26425 ( .A1(g25923), .A2(g9958), .ZN(g26425) );
AND2_X4 U_g26426 ( .A1(g5115), .A2(g25755), .ZN(g26426) );
AND2_X4 U_g26427 ( .A1(g5118), .A2(g25758), .ZN(g26427) );
AND2_X4 U_g26432 ( .A1(g5145), .A2(g25767), .ZN(g26432) );
AND2_X4 U_g26437 ( .A1(g5156), .A2(g25773), .ZN(g26437) );
AND2_X4 U_g26438 ( .A1(g5159), .A2(g25776), .ZN(g26438) );
AND2_X4 U_g26441 ( .A1(g5170), .A2(g25784), .ZN(g26441) );
AND2_X4 U_g26445 ( .A1(g5176), .A2(g25787), .ZN(g26445) );
AND2_X4 U_g26446 ( .A1(g5179), .A2(g25790), .ZN(g26446) );
AND2_X4 U_g26447 ( .A1(g5182), .A2(g25793), .ZN(g26447) );
AND2_X4 U_g26449 ( .A1(g5201), .A2(g25802), .ZN(g26449) );
AND2_X4 U_g26450 ( .A1(g5204), .A2(g25805), .ZN(g26450) );
AND2_X4 U_g26455 ( .A1(g5207), .A2(g25808), .ZN(g26455) );
AND2_X4 U_g26456 ( .A1(g5210), .A2(g25811), .ZN(g26456) );
AND2_X4 U_g26457 ( .A1(g5213), .A2(g25814), .ZN(g26457) );
AND2_X4 U_g26464 ( .A1(g5238), .A2(g25821), .ZN(g26464) );
AND2_X4 U_g26469 ( .A1(g5249), .A2(g25827), .ZN(g26469) );
AND2_X4 U_g26470 ( .A1(g5252), .A2(g25830), .ZN(g26470) );
AND2_X4 U_g26473 ( .A1(g5263), .A2(g25838), .ZN(g26473) );
AND2_X4 U_g26477 ( .A1(g5269), .A2(g25841), .ZN(g26477) );
AND2_X4 U_g26478 ( .A1(g5272), .A2(g25844), .ZN(g26478) );
AND2_X4 U_g26479 ( .A1(g5275), .A2(g25847), .ZN(g26479) );
AND2_X4 U_g26488 ( .A1(g5301), .A2(g25856), .ZN(g26488) );
AND2_X4 U_g26493 ( .A1(g5312), .A2(g25862), .ZN(g26493) );
AND2_X4 U_g26494 ( .A1(g5315), .A2(g25865), .ZN(g26494) );
AND2_X4 U_g26504 ( .A1(g5338), .A2(g25877), .ZN(g26504) );
AND2_X4 U_g26663 ( .A1(g25274), .A2(g21066), .ZN(g26663) );
AND2_X4 U_g26668 ( .A1(g25283), .A2(g21076), .ZN(g26668) );
AND2_X4 U_g26673 ( .A1(g12431), .A2(g25318), .ZN(g26673) );
AND2_X4 U_g26674 ( .A1(g25291), .A2(g21090), .ZN(g26674) );
AND2_X4 U_g26754 ( .A1(g14657), .A2(g26508), .ZN(g26754) );
AND2_X4 U_g26755 ( .A1(g26083), .A2(g22239), .ZN(g26755) );
AND2_X4 U_g26756 ( .A1(g26113), .A2(g22240), .ZN(g26756) );
AND3_X4 U_g26758 ( .A1(g16614), .A2(g26521), .A3(g13637), .ZN(g26758) );
AND2_X4 U_g26759 ( .A1(g26356), .A2(g19251), .ZN(g26759) );
AND2_X4 U_g26760 ( .A1(g26137), .A2(g22256), .ZN(g26760) );
AND2_X4 U_g26761 ( .A1(g26154), .A2(g22257), .ZN(g26761) );
AND2_X4 U_g26763 ( .A1(g14691), .A2(g26516), .ZN(g26763) );
AND3_X4 U_g26764 ( .A1(g16632), .A2(g26525), .A3(g13649), .ZN(g26764) );
AND2_X4 U_g26765 ( .A1(g26399), .A2(g19265), .ZN(g26765) );
AND2_X4 U_g26766 ( .A1(g14725), .A2(g26521), .ZN(g26766) );
AND2_X4 U_g26767 ( .A1(g26087), .A2(g22287), .ZN(g26767) );
AND2_X4 U_g26768 ( .A1(g26440), .A2(g19280), .ZN(g26768) );
AND2_X4 U_g26769 ( .A1(g14753), .A2(g26525), .ZN(g26769) );
AND2_X4 U_g26770 ( .A1(g26059), .A2(g19287), .ZN(g26770) );
AND3_X4 U_g26771 ( .A1(g24912), .A2(g26508), .A3(g13614), .ZN(g26771) );
AND2_X4 U_g26773 ( .A1(g26145), .A2(g22303), .ZN(g26773) );
AND2_X4 U_g26774 ( .A1(g26472), .A2(g19299), .ZN(g26774) );
AND2_X4 U_g26775 ( .A1(g26099), .A2(g22318), .ZN(g26775) );
AND2_X4 U_g26777 ( .A1(g26066), .A2(g19305), .ZN(g26777) );
AND3_X4 U_g26778 ( .A1(g24929), .A2(g26516), .A3(g13626), .ZN(g26778) );
AND2_X4 U_g26780 ( .A1(g26119), .A2(g16622), .ZN(g26780) );
AND2_X4 U_g26783 ( .A1(g26073), .A2(g19326), .ZN(g26783) );
AND3_X4 U_g26784 ( .A1(g24941), .A2(g26521), .A3(g13637), .ZN(g26784) );
AND2_X4 U_g26787 ( .A1(g26129), .A2(g16636), .ZN(g26787) );
AND2_X4 U_g26790 ( .A1(g26079), .A2(g19353), .ZN(g26790) );
AND3_X4 U_g26791 ( .A1(g24952), .A2(g26525), .A3(g13649), .ZN(g26791) );
AND2_X4 U_g26794 ( .A1(g26143), .A2(g16647), .ZN(g26794) );
AND2_X4 U_g26797 ( .A1(g26148), .A2(g16659), .ZN(g26797) );
AND2_X4 U_g26829 ( .A1(g5623), .A2(g26209), .ZN(g26829) );
AND2_X4 U_g26833 ( .A1(g5651), .A2(g26237), .ZN(g26833) );
AND2_X4 U_g26842 ( .A1(g5689), .A2(g26275), .ZN(g26842) );
AND2_X4 U_g26845 ( .A1(g5664), .A2(g26056), .ZN(g26845) );
AND2_X4 U_g26851 ( .A1(g5741), .A2(g26313), .ZN(g26851) );
AND2_X4 U_g26853 ( .A1(g5716), .A2(g26063), .ZN(g26853) );
AND2_X4 U_g26860 ( .A1(g5774), .A2(g26070), .ZN(g26860) );
AND2_X4 U_g26866 ( .A1(g5833), .A2(g26076), .ZN(g26866) );
AND2_X4 U_g26955 ( .A1(g6157), .A2(g26533), .ZN(g26955) );
AND2_X4 U_g26958 ( .A1(g6184), .A2(g26538), .ZN(g26958) );
AND2_X4 U_g26961 ( .A1(g13907), .A2(g26175), .ZN(g26961) );
AND2_X4 U_g26962 ( .A1(g6180), .A2(g26178), .ZN(g26962) );
AND2_X4 U_g26963 ( .A1(g6216), .A2(g26539), .ZN(g26963) );
AND2_X4 U_g26965 ( .A1(g23320), .A2(g26540), .ZN(g26965) );
AND2_X4 U_g26966 ( .A1(g13963), .A2(g26196), .ZN(g26966) );
AND2_X4 U_g26967 ( .A1(g6212), .A2(g26202), .ZN(g26967) );
AND2_X4 U_g26968 ( .A1(g6305), .A2(g26542), .ZN(g26968) );
AND2_X4 U_g26969 ( .A1(g23320), .A2(g26543), .ZN(g26969) );
AND2_X4 U_g26970 ( .A1(g21976), .A2(g26544), .ZN(g26970) );
AND2_X4 U_g26971 ( .A1(g23325), .A2(g26546), .ZN(g26971) );
AND2_X4 U_g26972 ( .A1(g14033), .A2(g26223), .ZN(g26972) );
AND2_X4 U_g26973 ( .A1(g6301), .A2(g26226), .ZN(g26973) );
AND2_X4 U_g26977 ( .A1(g23320), .A2(g26550), .ZN(g26977) );
AND2_X4 U_g26978 ( .A1(g21976), .A2(g26551), .ZN(g26978) );
AND2_X4 U_g26979 ( .A1(g23331), .A2(g26552), .ZN(g26979) );
AND2_X4 U_g26980 ( .A1(g23360), .A2(g26554), .ZN(g26980) );
AND2_X4 U_g26981 ( .A1(g23325), .A2(g26555), .ZN(g26981) );
AND2_X4 U_g26982 ( .A1(g21983), .A2(g26556), .ZN(g26982) );
AND2_X4 U_g26984 ( .A1(g23335), .A2(g26558), .ZN(g26984) );
AND2_X4 U_g26985 ( .A1(g14124), .A2(g26251), .ZN(g26985) );
AND2_X4 U_g26986 ( .A1(g6438), .A2(g26254), .ZN(g26986) );
AND2_X4 U_g26993 ( .A1(g21976), .A2(g26561), .ZN(g26993) );
AND2_X4 U_g26994 ( .A1(g23331), .A2(g26562), .ZN(g26994) );
AND2_X4 U_g26995 ( .A1(g21991), .A2(g26563), .ZN(g26995) );
AND2_X4 U_g26996 ( .A1(g23360), .A2(g26564), .ZN(g26996) );
AND2_X4 U_g26997 ( .A1(g22050), .A2(g26565), .ZN(g26997) );
AND2_X4 U_g26998 ( .A1(g23325), .A2(g26566), .ZN(g26998) );
AND2_X4 U_g26999 ( .A1(g21983), .A2(g26567), .ZN(g26999) );
AND2_X4 U_g27000 ( .A1(g23340), .A2(g26568), .ZN(g27000) );
AND2_X4 U_g27001 ( .A1(g23364), .A2(g26570), .ZN(g27001) );
AND2_X4 U_g27002 ( .A1(g23335), .A2(g26571), .ZN(g27002) );
AND2_X4 U_g27003 ( .A1(g21996), .A2(g26572), .ZN(g27003) );
AND2_X4 U_g27004 ( .A1(g23344), .A2(g26574), .ZN(g27004) );
AND2_X4 U_g27005 ( .A1(g23331), .A2(g26578), .ZN(g27005) );
AND2_X4 U_g27006 ( .A1(g21991), .A2(g26579), .ZN(g27006) );
AND2_X4 U_g27007 ( .A1(g23360), .A2(g26580), .ZN(g27007) );
AND2_X4 U_g27008 ( .A1(g22050), .A2(g26581), .ZN(g27008) );
AND2_X4 U_g27009 ( .A1(g23368), .A2(g26582), .ZN(g27009) );
AND2_X4 U_g27016 ( .A1(g21983), .A2(g26584), .ZN(g27016) );
AND2_X4 U_g27017 ( .A1(g23340), .A2(g26585), .ZN(g27017) );
AND2_X4 U_g27018 ( .A1(g22005), .A2(g26586), .ZN(g27018) );
AND2_X4 U_g27019 ( .A1(g23364), .A2(g26587), .ZN(g27019) );
AND2_X4 U_g27020 ( .A1(g22069), .A2(g26588), .ZN(g27020) );
AND2_X4 U_g27021 ( .A1(g23335), .A2(g26589), .ZN(g27021) );
AND2_X4 U_g27022 ( .A1(g21996), .A2(g26590), .ZN(g27022) );
AND2_X4 U_g27023 ( .A1(g23349), .A2(g26591), .ZN(g27023) );
AND2_X4 U_g27024 ( .A1(g23372), .A2(g26593), .ZN(g27024) );
AND2_X4 U_g27025 ( .A1(g23344), .A2(g26594), .ZN(g27025) );
AND2_X4 U_g27026 ( .A1(g22009), .A2(g26595), .ZN(g27026) );
AND2_X4 U_g27027 ( .A1(g21991), .A2(g26598), .ZN(g27027) );
AND2_X4 U_g27028 ( .A1(g22050), .A2(g26599), .ZN(g27028) );
AND2_X4 U_g27029 ( .A1(g23368), .A2(g26600), .ZN(g27029) );
AND2_X4 U_g27030 ( .A1(g22083), .A2(g26601), .ZN(g27030) );
AND2_X4 U_g27031 ( .A1(g23340), .A2(g26602), .ZN(g27031) );
AND2_X4 U_g27032 ( .A1(g22005), .A2(g26603), .ZN(g27032) );
AND2_X4 U_g27033 ( .A1(g23364), .A2(g26604), .ZN(g27033) );
AND2_X4 U_g27034 ( .A1(g22069), .A2(g26605), .ZN(g27034) );
AND2_X4 U_g27035 ( .A1(g23377), .A2(g26606), .ZN(g27035) );
AND2_X4 U_g27042 ( .A1(g21996), .A2(g26608), .ZN(g27042) );
AND2_X4 U_g27043 ( .A1(g23349), .A2(g26609), .ZN(g27043) );
AND2_X4 U_g27044 ( .A1(g22016), .A2(g26610), .ZN(g27044) );
AND2_X4 U_g27045 ( .A1(g23372), .A2(g26611), .ZN(g27045) );
AND2_X4 U_g27046 ( .A1(g22093), .A2(g26612), .ZN(g27046) );
AND2_X4 U_g27047 ( .A1(g23344), .A2(g26613), .ZN(g27047) );
AND2_X4 U_g27048 ( .A1(g22009), .A2(g26614), .ZN(g27048) );
AND2_X4 U_g27049 ( .A1(g23353), .A2(g26615), .ZN(g27049) );
AND2_X4 U_g27050 ( .A1(g23381), .A2(g26617), .ZN(g27050) );
AND2_X4 U_g27052 ( .A1(g4885), .A2(g26358), .ZN(g27052) );
AND2_X4 U_g27053 ( .A1(g23368), .A2(g26619), .ZN(g27053) );
AND2_X4 U_g27054 ( .A1(g22083), .A2(g26620), .ZN(g27054) );
AND2_X4 U_g27055 ( .A1(g22005), .A2(g26621), .ZN(g27055) );
AND2_X4 U_g27056 ( .A1(g22069), .A2(g26622), .ZN(g27056) );
AND2_X4 U_g27057 ( .A1(g23377), .A2(g26623), .ZN(g27057) );
AND2_X4 U_g27058 ( .A1(g22108), .A2(g26624), .ZN(g27058) );
AND2_X4 U_g27059 ( .A1(g23349), .A2(g26625), .ZN(g27059) );
AND2_X4 U_g27060 ( .A1(g22016), .A2(g26626), .ZN(g27060) );
AND2_X4 U_g27061 ( .A1(g23372), .A2(g26627), .ZN(g27061) );
AND2_X4 U_g27062 ( .A1(g22093), .A2(g26628), .ZN(g27062) );
AND2_X4 U_g27063 ( .A1(g23388), .A2(g26629), .ZN(g27063) );
AND2_X4 U_g27070 ( .A1(g22009), .A2(g26631), .ZN(g27070) );
AND2_X4 U_g27071 ( .A1(g23353), .A2(g26632), .ZN(g27071) );
AND2_X4 U_g27072 ( .A1(g22021), .A2(g26633), .ZN(g27072) );
AND2_X4 U_g27073 ( .A1(g23381), .A2(g26634), .ZN(g27073) );
AND2_X4 U_g27074 ( .A1(g22118), .A2(g26635), .ZN(g27074) );
AND2_X4 U_g27076 ( .A1(g5024), .A2(g26393), .ZN(g27076) );
AND2_X4 U_g27077 ( .A1(g22083), .A2(g26636), .ZN(g27077) );
AND2_X4 U_g27079 ( .A1(g5044), .A2(g26401), .ZN(g27079) );
AND2_X4 U_g27080 ( .A1(g23377), .A2(g26637), .ZN(g27080) );
AND2_X4 U_g27081 ( .A1(g22108), .A2(g26638), .ZN(g27081) );
AND2_X4 U_g27082 ( .A1(g22016), .A2(g26639), .ZN(g27082) );
AND2_X4 U_g27083 ( .A1(g22093), .A2(g26640), .ZN(g27083) );
AND2_X4 U_g27084 ( .A1(g23388), .A2(g26641), .ZN(g27084) );
AND2_X4 U_g27085 ( .A1(g22134), .A2(g26642), .ZN(g27085) );
AND2_X4 U_g27086 ( .A1(g23353), .A2(g26643), .ZN(g27086) );
AND2_X4 U_g27087 ( .A1(g22021), .A2(g26644), .ZN(g27087) );
AND2_X4 U_g27088 ( .A1(g23381), .A2(g26645), .ZN(g27088) );
AND2_X4 U_g27089 ( .A1(g22118), .A2(g26646), .ZN(g27089) );
AND2_X4 U_g27090 ( .A1(g23395), .A2(g26647), .ZN(g27090) );
AND2_X4 U_g27091 ( .A1(g5142), .A2(g26429), .ZN(g27091) );
AND2_X4 U_g27092 ( .A1(g5153), .A2(g26434), .ZN(g27092) );
AND2_X4 U_g27093 ( .A1(g22108), .A2(g26648), .ZN(g27093) );
AND2_X4 U_g27095 ( .A1(g5173), .A2(g26442), .ZN(g27095) );
AND2_X4 U_g27096 ( .A1(g23388), .A2(g26649), .ZN(g27096) );
AND2_X4 U_g27097 ( .A1(g22134), .A2(g26650), .ZN(g27097) );
AND2_X4 U_g27098 ( .A1(g22021), .A2(g26651), .ZN(g27098) );
AND2_X4 U_g27099 ( .A1(g22118), .A2(g26652), .ZN(g27099) );
AND2_X4 U_g27100 ( .A1(g23395), .A2(g26653), .ZN(g27100) );
AND2_X4 U_g27101 ( .A1(g22157), .A2(g26654), .ZN(g27101) );
AND2_X4 U_g27103 ( .A1(g5235), .A2(g26461), .ZN(g27103) );
AND2_X4 U_g27104 ( .A1(g5246), .A2(g26466), .ZN(g27104) );
AND2_X4 U_g27105 ( .A1(g22134), .A2(g26656), .ZN(g27105) );
AND2_X4 U_g27107 ( .A1(g5266), .A2(g26474), .ZN(g27107) );
AND2_X4 U_g27108 ( .A1(g23395), .A2(g26657), .ZN(g27108) );
AND2_X4 U_g27109 ( .A1(g22157), .A2(g26658), .ZN(g27109) );
AND2_X4 U_g27110 ( .A1(g5298), .A2(g26485), .ZN(g27110) );
AND2_X4 U_g27111 ( .A1(g5309), .A2(g26490), .ZN(g27111) );
AND2_X4 U_g27112 ( .A1(g22157), .A2(g26662), .ZN(g27112) );
AND2_X4 U_g27115 ( .A1(g5335), .A2(g26501), .ZN(g27115) );
AND2_X4 U_g27178 ( .A1(g26110), .A2(g22213), .ZN(g27178) );
AND3_X4 U_g27181 ( .A1(g16570), .A2(g26508), .A3(g13614), .ZN(g27181) );
AND2_X4 U_g27182 ( .A1(g26151), .A2(g22217), .ZN(g27182) );
AND2_X4 U_g27185 ( .A1(g26126), .A2(g22230), .ZN(g27185) );
AND3_X4 U_g27187 ( .A1(g16594), .A2(g26516), .A3(g13626), .ZN(g27187) );
AND2_X4 U_g27240 ( .A1(g26905), .A2(g22241), .ZN(g27240) );
AND2_X4 U_g27241 ( .A1(g10730), .A2(g26934), .ZN(g27241) );
AND2_X4 U_g27242 ( .A1(g26793), .A2(g8357), .ZN(g27242) );
AND2_X4 U_g27244 ( .A1(g26914), .A2(g22258), .ZN(g27244) );
AND2_X4 U_g27245 ( .A1(g26877), .A2(g22286), .ZN(g27245) );
AND2_X4 U_g27246 ( .A1(g26988), .A2(g16676), .ZN(g27246) );
AND2_X4 U_g27247 ( .A1(g27011), .A2(g16702), .ZN(g27247) );
AND2_X4 U_g27248 ( .A1(g27037), .A2(g16733), .ZN(g27248) );
AND2_X4 U_g27249 ( .A1(g27065), .A2(g16775), .ZN(g27249) );
AND2_X4 U_g27355 ( .A1(g61), .A2(g26837), .ZN(g27355) );
AND2_X4 U_g27356 ( .A1(g65), .A2(g26987), .ZN(g27356) );
AND2_X4 U_g27358 ( .A1(g749), .A2(g26846), .ZN(g27358) );
AND2_X4 U_g27359 ( .A1(g753), .A2(g27010), .ZN(g27359) );
AND2_X4 U_g27364 ( .A1(g1435), .A2(g26855), .ZN(g27364) );
AND2_X4 U_g27365 ( .A1(g1439), .A2(g27036), .ZN(g27365) );
AND2_X4 U_g27370 ( .A1(g27126), .A2(g8874), .ZN(g27370) );
AND2_X4 U_g27371 ( .A1(g2129), .A2(g26861), .ZN(g27371) );
AND2_X4 U_g27372 ( .A1(g2133), .A2(g27064), .ZN(g27372) );
AND2_X4 U_g27394 ( .A1(g17802), .A2(g27134), .ZN(g27394) );
AND2_X4 U_g27396 ( .A1(g692), .A2(g27135), .ZN(g27396) );
AND2_X4 U_g27407 ( .A1(g17914), .A2(g27136), .ZN(g27407) );
AND2_X4 U_g27409 ( .A1(g1378), .A2(g27137), .ZN(g27409) );
AND2_X4 U_g27425 ( .A1(g18025), .A2(g27138), .ZN(g27425) );
AND2_X4 U_g27427 ( .A1(g2072), .A2(g27139), .ZN(g27427) );
AND2_X4 U_g27446 ( .A1(g18142), .A2(g27141), .ZN(g27446) );
AND2_X4 U_g27448 ( .A1(g2766), .A2(g27142), .ZN(g27448) );
AND2_X4 U_g27495 ( .A1(g23945), .A2(g27146), .ZN(g27495) );
AND2_X4 U_g27509 ( .A1(g23945), .A2(g27148), .ZN(g27509) );
AND2_X4 U_g27516 ( .A1(g23974), .A2(g27151), .ZN(g27516) );
AND2_X4 U_g27530 ( .A1(g23945), .A2(g27153), .ZN(g27530) );
AND2_X4 U_g27534 ( .A1(g23974), .A2(g27155), .ZN(g27534) );
AND2_X4 U_g27541 ( .A1(g24004), .A2(g27159), .ZN(g27541) );
AND2_X4 U_g27552 ( .A1(g23974), .A2(g27162), .ZN(g27552) );
AND2_X4 U_g27554 ( .A1(g24004), .A2(g27164), .ZN(g27554) );
AND2_X4 U_g27561 ( .A1(g24038), .A2(g27167), .ZN(g27561) );
AND2_X4 U_g27568 ( .A1(g24004), .A2(g27172), .ZN(g27568) );
AND2_X4 U_g27570 ( .A1(g24038), .A2(g27173), .ZN(g27570) );
AND2_X4 U_g27578 ( .A1(g24038), .A2(g27177), .ZN(g27578) );
AND2_X4 U_g27656 ( .A1(g26796), .A2(g11004), .ZN(g27656) );
AND2_X4 U_g27657 ( .A1(g27114), .A2(g11051), .ZN(g27657) );
AND2_X4 U_g27659 ( .A1(g27132), .A2(g11114), .ZN(g27659) );
AND2_X4 U_g27660 ( .A1(g26835), .A2(g11117), .ZN(g27660) );
AND2_X4 U_g27661 ( .A1(g26841), .A2(g11173), .ZN(g27661) );
AND2_X4 U_g27666 ( .A1(g26849), .A2(g11243), .ZN(g27666) );
AND2_X4 U_g27671 ( .A1(g26885), .A2(g22212), .ZN(g27671) );
AND2_X4 U_g27673 ( .A1(g26854), .A2(g11312), .ZN(g27673) );
AND2_X4 U_g27679 ( .A1(g26782), .A2(g11386), .ZN(g27679) );
AND2_X4 U_g27680 ( .A1(g26983), .A2(g11392), .ZN(g27680) );
AND2_X4 U_g27681 ( .A1(g26788), .A2(g11456), .ZN(g27681) );
AND2_X4 U_g27719 ( .A1(g27496), .A2(g20649), .ZN(g27719) );
AND2_X4 U_g27720 ( .A1(g27481), .A2(g20652), .ZN(g27720) );
AND2_X4 U_g27721 ( .A1(g27579), .A2(g20655), .ZN(g27721) );
AND2_X4 U_g27723 ( .A1(g27464), .A2(g20679), .ZN(g27723) );
AND2_X4 U_g27725 ( .A1(g27532), .A2(g20704), .ZN(g27725) );
AND2_X4 U_g27726 ( .A1(g27531), .A2(g20732), .ZN(g27726) );
AND2_X4 U_g27727 ( .A1(g27414), .A2(g19301), .ZN(g27727) );
AND2_X4 U_g27728 ( .A1(g27564), .A2(g20766), .ZN(g27728) );
AND2_X4 U_g27729 ( .A1(g27435), .A2(g19322), .ZN(g27729) );
AND2_X4 U_g27730 ( .A1(g27454), .A2(g19349), .ZN(g27730) );
AND2_X4 U_g27731 ( .A1(g27470), .A2(g19383), .ZN(g27731) );
AND2_X4 U_g27732 ( .A1(g27492), .A2(g16758), .ZN(g27732) );
AND2_X4 U_g27733 ( .A1(g27513), .A2(g16785), .ZN(g27733) );
AND2_X4 U_g27734 ( .A1(g27538), .A2(g16814), .ZN(g27734) );
AND2_X4 U_g27737 ( .A1(g27558), .A2(g16832), .ZN(g27737) );
AND2_X4 U_g27770 ( .A1(g5642), .A2(g27449), .ZN(g27770) );
AND2_X4 U_g27772 ( .A1(g5680), .A2(g27465), .ZN(g27772) );
AND2_X4 U_g27773 ( .A1(g5732), .A2(g27484), .ZN(g27773) );
AND2_X4 U_g27774 ( .A1(g5702), .A2(g27361), .ZN(g27774) );
AND2_X4 U_g27775 ( .A1(g5790), .A2(g27506), .ZN(g27775) );
AND2_X4 U_g27779 ( .A1(g5760), .A2(g27367), .ZN(g27779) );
AND2_X4 U_g27783 ( .A1(g5819), .A2(g27373), .ZN(g27783) );
AND2_X4 U_g27790 ( .A1(g5875), .A2(g27376), .ZN(g27790) );
AND2_X4 U_g27904 ( .A1(g13873), .A2(g27387), .ZN(g27904) );
AND2_X4 U_g27908 ( .A1(g13886), .A2(g27391), .ZN(g27908) );
AND2_X4 U_g27909 ( .A1(g13895), .A2(g27397), .ZN(g27909) );
AND2_X4 U_g27913 ( .A1(g4017), .A2(g27401), .ZN(g27913) );
AND2_X4 U_g27914 ( .A1(g13927), .A2(g27404), .ZN(g27914) );
AND2_X4 U_g27915 ( .A1(g13936), .A2(g27410), .ZN(g27915) );
AND2_X4 U_g27922 ( .A1(g4112), .A2(g27416), .ZN(g27922) );
AND2_X4 U_g27923 ( .A1(g4144), .A2(g27419), .ZN(g27923) );
AND2_X4 U_g27924 ( .A1(g13983), .A2(g27422), .ZN(g27924) );
AND2_X4 U_g27926 ( .A1(g13992), .A2(g27428), .ZN(g27926) );
AND2_X4 U_g27931 ( .A1(g4221), .A2(g27432), .ZN(g27931) );
AND2_X4 U_g27935 ( .A1(g4251), .A2(g27437), .ZN(g27935) );
AND2_X4 U_g27936 ( .A1(g4283), .A2(g27440), .ZN(g27936) );
AND2_X4 U_g27938 ( .A1(g14053), .A2(g27443), .ZN(g27938) );
AND2_X4 U_g27945 ( .A1(g4376), .A2(g27451), .ZN(g27945) );
AND2_X4 U_g27949 ( .A1(g4406), .A2(g27456), .ZN(g27949) );
AND2_X4 U_g27951 ( .A1(g4438), .A2(g27459), .ZN(g27951) );
AND2_X4 U_g27963 ( .A1(g4545), .A2(g27467), .ZN(g27963) );
AND2_X4 U_g27968 ( .A1(g4575), .A2(g27472), .ZN(g27968) );
AND2_X4 U_g27970 ( .A1(g14238), .A2(g27475), .ZN(g27970) );
AND2_X4 U_g27984 ( .A1(g4721), .A2(g27486), .ZN(g27984) );
AND2_X4 U_g27985 ( .A1(g14342), .A2(g27489), .ZN(g27985) );
AND2_X4 U_g27991 ( .A1(g14360), .A2(g27498), .ZN(g27991) );
AND2_X4 U_g28008 ( .A1(g27590), .A2(g9770), .ZN(g28008) );
AND2_X4 U_g28009 ( .A1(g14454), .A2(g27510), .ZN(g28009) );
AND2_X4 U_g28015 ( .A1(g14472), .A2(g27518), .ZN(g28015) );
AND2_X4 U_g28027 ( .A1(g27590), .A2(g9895), .ZN(g28027) );
AND2_X4 U_g28028 ( .A1(g27595), .A2(g9898), .ZN(g28028) );
AND2_X4 U_g28035 ( .A1(g27599), .A2(g9916), .ZN(g28035) );
AND2_X4 U_g28036 ( .A1(g14541), .A2(g27535), .ZN(g28036) );
AND2_X4 U_g28042 ( .A1(g14559), .A2(g27543), .ZN(g28042) );
AND2_X4 U_g28050 ( .A1(g27590), .A2(g10018), .ZN(g28050) );
AND2_X4 U_g28051 ( .A1(g27595), .A2(g10021), .ZN(g28051) );
AND2_X4 U_g28057 ( .A1(g27599), .A2(g10049), .ZN(g28057) );
AND2_X4 U_g28058 ( .A1(g27604), .A2(g10052), .ZN(g28058) );
AND2_X4 U_g28065 ( .A1(g27608), .A2(g10070), .ZN(g28065) );
AND2_X4 U_g28066 ( .A1(g14596), .A2(g27555), .ZN(g28066) );
AND2_X4 U_g28073 ( .A1(g27595), .A2(g10109), .ZN(g28073) );
AND2_X4 U_g28079 ( .A1(g27599), .A2(g10127), .ZN(g28079) );
AND2_X4 U_g28080 ( .A1(g27604), .A2(g10130), .ZN(g28080) );
AND2_X4 U_g28086 ( .A1(g27608), .A2(g10158), .ZN(g28086) );
AND2_X4 U_g28087 ( .A1(g27613), .A2(g10161), .ZN(g28087) );
AND2_X4 U_g28094 ( .A1(g27617), .A2(g10179), .ZN(g28094) );
AND2_X4 U_g28098 ( .A1(g27604), .A2(g10214), .ZN(g28098) );
AND2_X4 U_g28104 ( .A1(g27608), .A2(g10232), .ZN(g28104) );
AND2_X4 U_g28105 ( .A1(g27613), .A2(g10235), .ZN(g28105) );
AND2_X4 U_g28111 ( .A1(g27617), .A2(g10263), .ZN(g28111) );
AND2_X4 U_g28112 ( .A1(g27622), .A2(g10266), .ZN(g28112) );
AND2_X4 U_g28116 ( .A1(g27613), .A2(g10316), .ZN(g28116) );
AND2_X4 U_g28122 ( .A1(g27617), .A2(g10334), .ZN(g28122) );
AND2_X4 U_g28123 ( .A1(g27622), .A2(g10337), .ZN(g28123) );
AND2_X4 U_g28127 ( .A1(g27622), .A2(g10409), .ZN(g28127) );
AND2_X4 U_g28171 ( .A1(g27349), .A2(g10898), .ZN(g28171) );
AND2_X4 U_g28176 ( .A1(g27349), .A2(g10940), .ZN(g28176) );
AND2_X4 U_g28188 ( .A1(g27349), .A2(g11008), .ZN(g28188) );
AND2_X4 U_g28193 ( .A1(g27573), .A2(g21914), .ZN(g28193) );
AND2_X4 U_g28319 ( .A1(g27855), .A2(g22246), .ZN(g28319) );
AND2_X4 U_g28320 ( .A1(g27854), .A2(g20637), .ZN(g28320) );
AND2_X4 U_g28322 ( .A1(g27937), .A2(g13868), .ZN(g28322) );
AND2_X4 U_g28323 ( .A1(g8580), .A2(g27838), .ZN(g28323) );
AND2_X4 U_g28324 ( .A1(g27810), .A2(g20659), .ZN(g28324) );
AND2_X4 U_g28326 ( .A1(g27865), .A2(g22274), .ZN(g28326) );
AND2_X4 U_g28327 ( .A1(g27900), .A2(g22275), .ZN(g28327) );
AND2_X4 U_g28329 ( .A1(g27823), .A2(g20708), .ZN(g28329) );
AND2_X4 U_g28330 ( .A1(g27864), .A2(g20711), .ZN(g28330) );
AND2_X4 U_g28331 ( .A1(g27802), .A2(g22307), .ZN(g28331) );
AND2_X4 U_g28332 ( .A1(g27883), .A2(g22331), .ZN(g28332) );
AND2_X4 U_g28333 ( .A1(g27882), .A2(g20772), .ZN(g28333) );
AND2_X4 U_g28334 ( .A1(g27842), .A2(g20793), .ZN(g28334) );
AND2_X4 U_g28335 ( .A1(g27814), .A2(g22343), .ZN(g28335) );
AND2_X4 U_g28336 ( .A1(g27896), .A2(g20810), .ZN(g28336) );
AND2_X4 U_g28337 ( .A1(g28002), .A2(g19448), .ZN(g28337) );
AND2_X4 U_g28338 ( .A1(g28029), .A2(g19475), .ZN(g28338) );
AND2_X4 U_g28339 ( .A1(g28059), .A2(g19498), .ZN(g28339) );
AND2_X4 U_g28340 ( .A1(g28088), .A2(g19519), .ZN(g28340) );
AND2_X4 U_g28373 ( .A1(g56), .A2(g27969), .ZN(g28373) );
AND2_X4 U_g28376 ( .A1(g744), .A2(g27990), .ZN(g28376) );
AND2_X4 U_g28378 ( .A1(g52), .A2(g27776), .ZN(g28378) );
AND3_X4 U_g28379 ( .A1(g27868), .A2(g19390), .A3(g19369), .ZN(g28379) );
AND2_X4 U_g28380 ( .A1(g1430), .A2(g28014), .ZN(g28380) );
AND2_X4 U_g28381 ( .A1(g28157), .A2(g9815), .ZN(g28381) );
AND2_X4 U_g28383 ( .A1(g740), .A2(g27780), .ZN(g28383) );
AND2_X4 U_g28385 ( .A1(g2124), .A2(g28041), .ZN(g28385) );
AND2_X4 U_g28387 ( .A1(g1426), .A2(g27787), .ZN(g28387) );
AND2_X4 U_g28389 ( .A1(g2120), .A2(g27794), .ZN(g28389) );
AND2_X4 U_g28396 ( .A1(g7754), .A2(g27806), .ZN(g28396) );
AND2_X4 U_g28398 ( .A1(g7769), .A2(g27817), .ZN(g28398) );
AND2_X4 U_g28399 ( .A1(g7776), .A2(g27820), .ZN(g28399) );
AND2_X4 U_g28401 ( .A1(g7782), .A2(g27831), .ZN(g28401) );
AND2_X4 U_g28402 ( .A1(g7785), .A2(g27839), .ZN(g28402) );
AND2_X4 U_g28404 ( .A1(g7792), .A2(g27843), .ZN(g28404) );
AND2_X4 U_g28405 ( .A1(g7796), .A2(g27847), .ZN(g28405) );
AND2_X4 U_g28407 ( .A1(g7799), .A2(g27858), .ZN(g28407) );
AND2_X4 U_g28408 ( .A1(g7806), .A2(g27861), .ZN(g28408) );
AND2_X4 U_g28411 ( .A1(g7809), .A2(g27872), .ZN(g28411) );
AND2_X4 U_g28412 ( .A1(g7812), .A2(g27879), .ZN(g28412) );
AND2_X4 U_g28416 ( .A1(g7823), .A2(g27889), .ZN(g28416) );
AND2_X4 U_g28422 ( .A1(g17640), .A2(g28150), .ZN(g28422) );
AND2_X4 U_g28423 ( .A1(g17724), .A2(g28152), .ZN(g28423) );
AND2_X4 U_g28424 ( .A1(g17741), .A2(g28153), .ZN(g28424) );
AND2_X4 U_g28426 ( .A1(g28128), .A2(g9170), .ZN(g28426) );
AND2_X4 U_g28427 ( .A1(g26092), .A2(g28154), .ZN(g28427) );
AND2_X4 U_g28428 ( .A1(g17825), .A2(g28155), .ZN(g28428) );
AND2_X4 U_g28429 ( .A1(g17842), .A2(g28156), .ZN(g28429) );
AND2_X4 U_g28430 ( .A1(g28128), .A2(g9196), .ZN(g28430) );
AND2_X4 U_g28431 ( .A1(g26092), .A2(g28158), .ZN(g28431) );
AND2_X4 U_g28433 ( .A1(g28133), .A2(g9212), .ZN(g28433) );
AND2_X4 U_g28434 ( .A1(g26114), .A2(g28159), .ZN(g28434) );
AND2_X4 U_g28435 ( .A1(g17937), .A2(g28160), .ZN(g28435) );
AND2_X4 U_g28436 ( .A1(g17954), .A2(g28161), .ZN(g28436) );
AND2_X4 U_g28438 ( .A1(g17882), .A2(g27919), .ZN(g28438) );
AND2_X4 U_g28439 ( .A1(g28128), .A2(g9242), .ZN(g28439) );
AND2_X4 U_g28440 ( .A1(g26092), .A2(g28162), .ZN(g28440) );
AND2_X4 U_g28441 ( .A1(g28133), .A2(g9257), .ZN(g28441) );
AND2_X4 U_g28442 ( .A1(g26114), .A2(g28163), .ZN(g28442) );
AND2_X4 U_g28444 ( .A1(g28137), .A2(g9273), .ZN(g28444) );
AND2_X4 U_g28445 ( .A1(g26121), .A2(g28164), .ZN(g28445) );
AND2_X4 U_g28446 ( .A1(g18048), .A2(g28165), .ZN(g28446) );
AND2_X4 U_g28448 ( .A1(g17974), .A2(g27928), .ZN(g28448) );
AND2_X4 U_g28450 ( .A1(g17993), .A2(g27932), .ZN(g28450) );
AND2_X4 U_g28451 ( .A1(g28133), .A2(g9320), .ZN(g28451) );
AND2_X4 U_g28452 ( .A1(g26114), .A2(g28166), .ZN(g28452) );
AND2_X4 U_g28453 ( .A1(g28137), .A2(g9335), .ZN(g28453) );
AND2_X4 U_g28454 ( .A1(g26121), .A2(g28167), .ZN(g28454) );
AND2_X4 U_g28456 ( .A1(g28141), .A2(g9351), .ZN(g28456) );
AND2_X4 U_g28457 ( .A1(g26131), .A2(g28168), .ZN(g28457) );
AND2_X4 U_g28459 ( .A1(g18074), .A2(g27939), .ZN(g28459) );
AND2_X4 U_g28460 ( .A1(g18091), .A2(g27942), .ZN(g28460) );
AND2_X4 U_g28462 ( .A1(g18110), .A2(g27946), .ZN(g28462) );
AND2_X4 U_g28463 ( .A1(g28137), .A2(g9401), .ZN(g28463) );
AND2_X4 U_g28464 ( .A1(g26121), .A2(g28169), .ZN(g28464) );
AND2_X4 U_g28465 ( .A1(g28141), .A2(g9416), .ZN(g28465) );
AND2_X4 U_g28466 ( .A1(g26131), .A2(g28170), .ZN(g28466) );
AND2_X4 U_g28468 ( .A1(g18265), .A2(g28172), .ZN(g28468) );
AND2_X4 U_g28469 ( .A1(g18179), .A2(g27952), .ZN(g28469) );
AND2_X4 U_g28471 ( .A1(g18190), .A2(g27956), .ZN(g28471) );
AND2_X4 U_g28472 ( .A1(g18207), .A2(g27959), .ZN(g28472) );
AND2_X4 U_g28474 ( .A1(g18226), .A2(g27965), .ZN(g28474) );
AND2_X4 U_g28475 ( .A1(g28141), .A2(g9498), .ZN(g28475) );
AND2_X4 U_g28476 ( .A1(g26131), .A2(g28173), .ZN(g28476) );
AND2_X4 U_g28477 ( .A1(g18341), .A2(g28174), .ZN(g28477) );
AND2_X4 U_g28478 ( .A1(g18358), .A2(g28175), .ZN(g28478) );
AND2_X4 U_g28479 ( .A1(g18286), .A2(g27973), .ZN(g28479) );
AND2_X4 U_g28480 ( .A1(g18297), .A2(g27977), .ZN(g28480) );
AND2_X4 U_g28481 ( .A1(g18314), .A2(g27981), .ZN(g28481) );
AND2_X4 U_g28484 ( .A1(g18436), .A2(g28177), .ZN(g28484) );
AND2_X4 U_g28485 ( .A1(g18453), .A2(g28178), .ZN(g28485) );
AND2_X4 U_g28486 ( .A1(g18379), .A2(g27994), .ZN(g28486) );
AND2_X4 U_g28487 ( .A1(g18390), .A2(g27999), .ZN(g28487) );
AND2_X4 U_g28492 ( .A1(g18509), .A2(g28186), .ZN(g28492) );
AND2_X4 U_g28493 ( .A1(g18526), .A2(g28187), .ZN(g28493) );
AND2_X4 U_g28494 ( .A1(g18474), .A2(g28018), .ZN(g28494) );
AND2_X4 U_g28497 ( .A1(g18573), .A2(g28190), .ZN(g28497) );
AND2_X4 U_g28657 ( .A1(g27925), .A2(g13700), .ZN(g28657) );
AND2_X4 U_g28659 ( .A1(g27917), .A2(g13736), .ZN(g28659) );
AND2_X4 U_g28660 ( .A1(g27916), .A2(g11911), .ZN(g28660) );
AND2_X4 U_g28662 ( .A1(g27911), .A2(g11951), .ZN(g28662) );
AND2_X4 U_g28663 ( .A1(g27906), .A2(g11997), .ZN(g28663) );
AND2_X4 U_g28664 ( .A1(g27997), .A2(g12055), .ZN(g28664) );
AND2_X4 U_g28665 ( .A1(g27827), .A2(g22222), .ZN(g28665) );
AND2_X4 U_g28666 ( .A1(g27980), .A2(g12106), .ZN(g28666) );
AND2_X4 U_g28667 ( .A1(g27964), .A2(g13852), .ZN(g28667) );
AND2_X4 U_g28669 ( .A1(g27897), .A2(g22233), .ZN(g28669) );
AND2_X4 U_g28670 ( .A1(g27798), .A2(g21935), .ZN(g28670) );
AND2_X4 U_g28671 ( .A1(g27962), .A2(g12161), .ZN(g28671) );
AND2_X4 U_g28672 ( .A1(g27950), .A2(g13859), .ZN(g28672) );
AND2_X4 U_g28707 ( .A1(g12436), .A2(g28379), .ZN(g28707) );
AND2_X4 U_g28708 ( .A1(g28392), .A2(g22260), .ZN(g28708) );
AND2_X4 U_g28709 ( .A1(g28400), .A2(g22261), .ZN(g28709) );
AND2_X4 U_g28710 ( .A1(g28403), .A2(g22262), .ZN(g28710) );
AND2_X4 U_g28711 ( .A1(g10749), .A2(g28415), .ZN(g28711) );
AND2_X4 U_g28712 ( .A1(g28406), .A2(g22276), .ZN(g28712) );
AND2_X4 U_g28713 ( .A1(g28410), .A2(g22290), .ZN(g28713) );
AND2_X4 U_g28714 ( .A1(g28394), .A2(g22306), .ZN(g28714) );
AND2_X4 U_g28715 ( .A1(g28414), .A2(g22332), .ZN(g28715) );
AND2_X4 U_g28716 ( .A1(g28449), .A2(g19319), .ZN(g28716) );
AND2_X4 U_g28717 ( .A1(g28461), .A2(g19346), .ZN(g28717) );
AND2_X4 U_g28718 ( .A1(g28473), .A2(g19380), .ZN(g28718) );
AND2_X4 U_g28719 ( .A1(g28482), .A2(g19412), .ZN(g28719) );
AND2_X4 U_g28722 ( .A1(g28523), .A2(g16694), .ZN(g28722) );
AND2_X4 U_g28724 ( .A1(g28551), .A2(g16725), .ZN(g28724) );
AND2_X4 U_g28726 ( .A1(g28578), .A2(g16767), .ZN(g28726) );
AND2_X4 U_g28729 ( .A1(g28606), .A2(g16794), .ZN(g28729) );
AND2_X4 U_g28834 ( .A1(g5751), .A2(g28483), .ZN(g28834) );
AND2_X4 U_g28836 ( .A1(g5810), .A2(g28491), .ZN(g28836) );
AND2_X4 U_g28838 ( .A1(g5866), .A2(g28496), .ZN(g28838) );
AND2_X4 U_g28840 ( .A1(g5913), .A2(g28500), .ZN(g28840) );
AND2_X4 U_g28841 ( .A1(g27834), .A2(g28554), .ZN(g28841) );
AND2_X4 U_g28843 ( .A1(g27834), .A2(g28581), .ZN(g28843) );
AND2_X4 U_g28844 ( .A1(g27850), .A2(g28582), .ZN(g28844) );
AND2_X4 U_g28846 ( .A1(g27834), .A2(g28608), .ZN(g28846) );
AND2_X4 U_g28847 ( .A1(g27850), .A2(g28609), .ZN(g28847) );
AND2_X4 U_g28848 ( .A1(g27875), .A2(g28610), .ZN(g28848) );
AND2_X4 U_g28849 ( .A1(g27850), .A2(g28616), .ZN(g28849) );
AND2_X4 U_g28850 ( .A1(g27875), .A2(g28617), .ZN(g28850) );
AND2_X4 U_g28851 ( .A1(g27892), .A2(g28618), .ZN(g28851) );
AND2_X4 U_g28852 ( .A1(g27875), .A2(g28623), .ZN(g28852) );
AND2_X4 U_g28853 ( .A1(g27892), .A2(g28624), .ZN(g28853) );
AND2_X4 U_g28854 ( .A1(g27892), .A2(g28629), .ZN(g28854) );
AND2_X4 U_g28880 ( .A1(g13946), .A2(g28639), .ZN(g28880) );
AND2_X4 U_g28881 ( .A1(g28612), .A2(g9199), .ZN(g28881) );
AND2_X4 U_g28892 ( .A1(g14001), .A2(g28640), .ZN(g28892) );
AND2_X4 U_g28893 ( .A1(g28612), .A2(g9245), .ZN(g28893) );
AND2_X4 U_g28897 ( .A1(g14016), .A2(g28641), .ZN(g28897) );
AND2_X4 U_g28898 ( .A1(g28619), .A2(g9260), .ZN(g28898) );
AND2_X4 U_g28909 ( .A1(g14062), .A2(g28642), .ZN(g28909) );
AND2_X4 U_g28910 ( .A1(g28612), .A2(g9303), .ZN(g28910) );
AND2_X4 U_g28914 ( .A1(g14092), .A2(g28643), .ZN(g28914) );
AND2_X4 U_g28915 ( .A1(g28619), .A2(g9323), .ZN(g28915) );
AND2_X4 U_g28919 ( .A1(g14107), .A2(g28644), .ZN(g28919) );
AND2_X4 U_g28923 ( .A1(g28625), .A2(g9338), .ZN(g28923) );
AND2_X4 U_g28931 ( .A1(g14153), .A2(g28645), .ZN(g28931) );
AND2_X4 U_g28935 ( .A1(g14177), .A2(g28646), .ZN(g28935) );
AND2_X4 U_g28936 ( .A1(g28619), .A2(g9384), .ZN(g28936) );
AND2_X4 U_g28940 ( .A1(g14207), .A2(g28647), .ZN(g28940) );
AND2_X4 U_g28944 ( .A1(g28625), .A2(g9404), .ZN(g28944) );
AND2_X4 U_g28948 ( .A1(g14222), .A2(g28648), .ZN(g28948) );
AND2_X4 U_g28949 ( .A1(g28630), .A2(g9419), .ZN(g28949) );
AND2_X4 U_g28958 ( .A1(g14268), .A2(g28649), .ZN(g28958) );
AND2_X4 U_g28962 ( .A1(g14292), .A2(g28650), .ZN(g28962) );
AND2_X4 U_g28966 ( .A1(g28625), .A2(g9481), .ZN(g28966) );
AND2_X4 U_g28970 ( .A1(g14322), .A2(g28651), .ZN(g28970) );
AND2_X4 U_g28971 ( .A1(g28630), .A2(g9501), .ZN(g28971) );
AND2_X4 U_g28986 ( .A1(g14390), .A2(g28652), .ZN(g28986) );
AND2_X4 U_g28996 ( .A1(g14414), .A2(g28653), .ZN(g28996) );
AND2_X4 U_g28997 ( .A1(g28630), .A2(g9623), .ZN(g28997) );
AND2_X4 U_g29022 ( .A1(g14502), .A2(g28655), .ZN(g29022) );
AND2_X4 U_g29130 ( .A1(g28397), .A2(g22221), .ZN(g29130) );
AND2_X4 U_g29174 ( .A1(g29031), .A2(g20684), .ZN(g29174) );
AND2_X4 U_g29175 ( .A1(g29009), .A2(g20687), .ZN(g29175) );
AND2_X4 U_g29176 ( .A1(g29097), .A2(g20690), .ZN(g29176) );
AND2_X4 U_g29180 ( .A1(g28982), .A2(g20714), .ZN(g29180) );
AND2_X4 U_g29183 ( .A1(g29064), .A2(g20739), .ZN(g29183) );
AND2_X4 U_g29186 ( .A1(g29063), .A2(g20769), .ZN(g29186) );
AND2_X4 U_g29188 ( .A1(g29083), .A2(g20796), .ZN(g29188) );
AND2_X4 U_g29196 ( .A1(g15022), .A2(g28741), .ZN(g29196) );
AND2_X4 U_g29200 ( .A1(g15096), .A2(g28751), .ZN(g29200) );
AND2_X4 U_g29203 ( .A1(g15118), .A2(g28755), .ZN(g29203) );
AND2_X4 U_g29208 ( .A1(g15188), .A2(g28764), .ZN(g29208) );
AND2_X4 U_g29211 ( .A1(g15210), .A2(g28768), .ZN(g29211) );
AND2_X4 U_g29217 ( .A1(g15274), .A2(g28775), .ZN(g29217) );
AND2_X4 U_g29220 ( .A1(g15296), .A2(g28779), .ZN(g29220) );
AND2_X4 U_g29225 ( .A1(g15366), .A2(g28785), .ZN(g29225) );
AND2_X4 U_g29229 ( .A1(g9293), .A2(g28791), .ZN(g29229) );
AND2_X4 U_g29232 ( .A1(g9356), .A2(g28796), .ZN(g29232) );
AND2_X4 U_g29233 ( .A1(g9374), .A2(g28799), .ZN(g29233) );
AND2_X4 U_g29234 ( .A1(g9427), .A2(g28804), .ZN(g29234) );
AND2_X4 U_g29235 ( .A1(g9453), .A2(g28807), .ZN(g29235) );
AND2_X4 U_g29236 ( .A1(g9471), .A2(g28810), .ZN(g29236) );
AND2_X4 U_g29238 ( .A1(g9569), .A2(g28814), .ZN(g29238) );
AND2_X4 U_g29239 ( .A1(g9595), .A2(g28817), .ZN(g29239) );
AND2_X4 U_g29240 ( .A1(g9613), .A2(g28820), .ZN(g29240) );
AND2_X4 U_g29241 ( .A1(g9711), .A2(g28823), .ZN(g29241) );
AND2_X4 U_g29242 ( .A1(g9737), .A2(g28826), .ZN(g29242) );
AND2_X4 U_g29243 ( .A1(g9857), .A2(g28829), .ZN(g29243) );
AND2_X4 U_g29248 ( .A1(g28855), .A2(g8836), .ZN(g29248) );
AND2_X4 U_g29251 ( .A1(g28855), .A2(g8856), .ZN(g29251) );
AND2_X4 U_g29252 ( .A1(g28859), .A2(g8863), .ZN(g29252) );
AND2_X4 U_g29255 ( .A1(g28855), .A2(g8885), .ZN(g29255) );
AND2_X4 U_g29256 ( .A1(g28859), .A2(g8894), .ZN(g29256) );
AND2_X4 U_g29257 ( .A1(g28863), .A2(g8901), .ZN(g29257) );
AND2_X4 U_g29259 ( .A1(g28859), .A2(g8925), .ZN(g29259) );
AND2_X4 U_g29260 ( .A1(g28863), .A2(g8934), .ZN(g29260) );
AND2_X4 U_g29261 ( .A1(g28867), .A2(g8941), .ZN(g29261) );
AND2_X4 U_g29262 ( .A1(g28863), .A2(g8965), .ZN(g29262) );
AND2_X4 U_g29263 ( .A1(g28867), .A2(g8974), .ZN(g29263) );
AND2_X4 U_g29264 ( .A1(g28867), .A2(g8997), .ZN(g29264) );
AND2_X4 U_g29284 ( .A1(g29001), .A2(g28871), .ZN(g29284) );
AND2_X4 U_g29289 ( .A1(g29030), .A2(g28883), .ZN(g29289) );
AND2_X4 U_g29294 ( .A1(g29053), .A2(g28900), .ZN(g29294) );
AND2_X4 U_g29300 ( .A1(g29072), .A2(g28925), .ZN(g29300) );
AND2_X4 U_g29302 ( .A1(g29026), .A2(g28928), .ZN(g29302) );
AND2_X4 U_g29310 ( .A1(g28978), .A2(g28951), .ZN(g29310) );
AND2_X4 U_g29312 ( .A1(g29049), .A2(g28955), .ZN(g29312) );
AND2_X4 U_g29320 ( .A1(g29088), .A2(g28972), .ZN(g29320) );
AND2_X4 U_g29321 ( .A1(g29008), .A2(g28979), .ZN(g29321) );
AND2_X4 U_g29323 ( .A1(g29068), .A2(g28983), .ZN(g29323) );
AND2_X4 U_g29329 ( .A1(g29096), .A2(g29002), .ZN(g29329) );
AND2_X4 U_g29330 ( .A1(g29038), .A2(g29010), .ZN(g29330) );
AND2_X4 U_g29332 ( .A1(g29080), .A2(g29019), .ZN(g29332) );
AND2_X4 U_g29336 ( .A1(g29045), .A2(g29023), .ZN(g29336) );
AND2_X4 U_g29337 ( .A1(g29103), .A2(g29032), .ZN(g29337) );
AND2_X4 U_g29338 ( .A1(g29060), .A2(g29042), .ZN(g29338) );
AND2_X4 U_g29341 ( .A1(g29062), .A2(g29046), .ZN(g29341) );
AND2_X4 U_g29342 ( .A1(g29107), .A2(g29054), .ZN(g29342) );
AND2_X4 U_g29344 ( .A1(g29076), .A2(g29065), .ZN(g29344) );
AND2_X4 U_g29346 ( .A1(g29087), .A2(g29077), .ZN(g29346) );
AND2_X4 U_g29411 ( .A1(g29090), .A2(g21932), .ZN(g29411) );
AND2_X4 U_g29464 ( .A1(g29190), .A2(g8375), .ZN(g29464) );
AND2_X4 U_g29465 ( .A1(g29191), .A2(g8424), .ZN(g29465) );
AND2_X4 U_g29466 ( .A1(g8587), .A2(g29265), .ZN(g29466) );
AND2_X4 U_g29467 ( .A1(g29340), .A2(g19467), .ZN(g29467) );
AND2_X4 U_g29468 ( .A1(g29343), .A2(g19490), .ZN(g29468) );
AND2_X4 U_g29469 ( .A1(g29345), .A2(g19511), .ZN(g29469) );
AND2_X4 U_g29470 ( .A1(g29347), .A2(g19530), .ZN(g29470) );
AND2_X4 U_g29471 ( .A1(g21461), .A2(g29266), .ZN(g29471) );
AND2_X4 U_g29472 ( .A1(g21461), .A2(g29268), .ZN(g29472) );
AND2_X4 U_g29473 ( .A1(g21508), .A2(g29269), .ZN(g29473) );
AND2_X4 U_g29474 ( .A1(g21508), .A2(g29271), .ZN(g29474) );
AND2_X4 U_g29475 ( .A1(g21544), .A2(g29272), .ZN(g29475) );
AND2_X4 U_g29476 ( .A1(g21544), .A2(g29274), .ZN(g29476) );
AND2_X4 U_g29477 ( .A1(g21580), .A2(g29275), .ZN(g29477) );
AND2_X4 U_g29478 ( .A1(g21580), .A2(g29277), .ZN(g29478) );
AND2_X4 U_g29479 ( .A1(g21461), .A2(g29280), .ZN(g29479) );
AND2_X4 U_g29480 ( .A1(g21461), .A2(g29282), .ZN(g29480) );
AND2_X4 U_g29481 ( .A1(g21508), .A2(g29283), .ZN(g29481) );
AND2_X4 U_g29482 ( .A1(g21461), .A2(g29285), .ZN(g29482) );
AND2_X4 U_g29483 ( .A1(g21508), .A2(g29286), .ZN(g29483) );
AND2_X4 U_g29484 ( .A1(g21544), .A2(g29287), .ZN(g29484) );
AND2_X4 U_g29485 ( .A1(g21508), .A2(g29290), .ZN(g29485) );
AND2_X4 U_g29486 ( .A1(g21544), .A2(g29291), .ZN(g29486) );
AND2_X4 U_g29487 ( .A1(g21580), .A2(g29292), .ZN(g29487) );
AND2_X4 U_g29488 ( .A1(g21544), .A2(g29295), .ZN(g29488) );
AND2_X4 U_g29489 ( .A1(g21580), .A2(g29296), .ZN(g29489) );
AND2_X4 U_g29490 ( .A1(g21580), .A2(g29301), .ZN(g29490) );
AND2_X4 U_g29502 ( .A1(g29350), .A2(g8912), .ZN(g29502) );
AND2_X4 U_g29518 ( .A1(g28728), .A2(g29360), .ZN(g29518) );
AND2_X4 U_g29520 ( .A1(g28731), .A2(g29361), .ZN(g29520) );
AND2_X4 U_g29521 ( .A1(g28733), .A2(g29362), .ZN(g29521) );
AND2_X4 U_g29522 ( .A1(g27735), .A2(g29363), .ZN(g29522) );
AND2_X4 U_g29523 ( .A1(g28737), .A2(g29364), .ZN(g29523) );
AND2_X4 U_g29524 ( .A1(g28739), .A2(g29365), .ZN(g29524) );
AND2_X4 U_g29525 ( .A1(g29195), .A2(g29366), .ZN(g29525) );
AND2_X4 U_g29526 ( .A1(g27741), .A2(g29367), .ZN(g29526) );
AND2_X4 U_g29527 ( .A1(g28748), .A2(g29368), .ZN(g29527) );
AND2_X4 U_g29528 ( .A1(g28750), .A2(g29369), .ZN(g29528) );
AND2_X4 U_g29529 ( .A1(g29199), .A2(g29370), .ZN(g29529) );
AND2_X4 U_g29531 ( .A1(g29202), .A2(g29371), .ZN(g29531) );
AND2_X4 U_g29532 ( .A1(g27746), .A2(g29372), .ZN(g29532) );
AND2_X4 U_g29533 ( .A1(g28762), .A2(g29373), .ZN(g29533) );
AND2_X4 U_g29534 ( .A1(g29206), .A2(g29374), .ZN(g29534) );
AND2_X4 U_g29536 ( .A1(g29207), .A2(g29375), .ZN(g29536) );
AND2_X4 U_g29538 ( .A1(g29210), .A2(g29376), .ZN(g29538) );
AND2_X4 U_g29539 ( .A1(g27754), .A2(g29377), .ZN(g29539) );
AND2_X4 U_g29540 ( .A1(g26041), .A2(g29378), .ZN(g29540) );
AND2_X4 U_g29541 ( .A1(g29214), .A2(g29379), .ZN(g29541) );
AND2_X4 U_g29543 ( .A1(g29215), .A2(g29380), .ZN(g29543) );
AND2_X4 U_g29545 ( .A1(g29216), .A2(g29381), .ZN(g29545) );
AND2_X4 U_g29547 ( .A1(g29219), .A2(g29382), .ZN(g29547) );
AND2_X4 U_g29548 ( .A1(g28784), .A2(g29383), .ZN(g29548) );
AND2_X4 U_g29549 ( .A1(g26043), .A2(g29384), .ZN(g29549) );
AND2_X4 U_g29550 ( .A1(g29222), .A2(g29385), .ZN(g29550) );
AND2_X4 U_g29553 ( .A1(g29223), .A2(g29386), .ZN(g29553) );
AND2_X4 U_g29555 ( .A1(g29224), .A2(g29387), .ZN(g29555) );
AND2_X4 U_g29557 ( .A1(g28789), .A2(g29388), .ZN(g29557) );
AND2_X4 U_g29558 ( .A1(g28790), .A2(g29389), .ZN(g29558) );
AND2_X4 U_g29559 ( .A1(g26045), .A2(g29390), .ZN(g29559) );
AND2_X4 U_g29560 ( .A1(g29227), .A2(g29391), .ZN(g29560) );
AND2_X4 U_g29562 ( .A1(g29228), .A2(g29392), .ZN(g29562) );
AND2_X4 U_g29564 ( .A1(g28794), .A2(g29393), .ZN(g29564) );
AND2_X4 U_g29565 ( .A1(g28795), .A2(g29394), .ZN(g29565) );
AND2_X4 U_g29566 ( .A1(g26047), .A2(g29395), .ZN(g29566) );
AND2_X4 U_g29567 ( .A1(g29231), .A2(g29396), .ZN(g29567) );
AND2_X4 U_g29572 ( .A1(g28802), .A2(g29397), .ZN(g29572) );
AND2_X4 U_g29573 ( .A1(g28803), .A2(g29398), .ZN(g29573) );
AND2_X4 U_g29575 ( .A1(g28813), .A2(g29402), .ZN(g29575) );
AND2_X4 U_g29607 ( .A1(g29193), .A2(g11056), .ZN(g29607) );
AND2_X4 U_g29610 ( .A1(g29349), .A2(g11123), .ZN(g29610) );
AND2_X4 U_g29614 ( .A1(g29359), .A2(g11182), .ZN(g29614) );
AND2_X4 U_g29615 ( .A1(g29245), .A2(g11185), .ZN(g29615) );
AND2_X4 U_g29619 ( .A1(g29247), .A2(g11259), .ZN(g29619) );
AND2_X4 U_g29622 ( .A1(g29250), .A2(g11327), .ZN(g29622) );
AND2_X4 U_g29624 ( .A1(g29254), .A2(g11407), .ZN(g29624) );
AND2_X4 U_g29625 ( .A1(g29189), .A2(g11472), .ZN(g29625) );
AND2_X4 U_g29626 ( .A1(g29318), .A2(g11478), .ZN(g29626) );
AND2_X4 U_g29790 ( .A1(g29491), .A2(g10918), .ZN(g29790) );
AND2_X4 U_g29792 ( .A1(g29491), .A2(g10977), .ZN(g29792) );
AND2_X4 U_g29793 ( .A1(g29491), .A2(g11063), .ZN(g29793) );
AND2_X4 U_g29810 ( .A1(g29748), .A2(g22248), .ZN(g29810) );
AND2_X4 U_g29811 ( .A1(g29703), .A2(g20644), .ZN(g29811) );
AND2_X4 U_g29812 ( .A1(g29762), .A2(g12223), .ZN(g29812) );
AND2_X4 U_g29813 ( .A1(g29760), .A2(g13869), .ZN(g29813) );
AND2_X4 U_g29814 ( .A1(g29728), .A2(g22266), .ZN(g29814) );
AND2_X4 U_g29815 ( .A1(g29727), .A2(g20662), .ZN(g29815) );
AND2_X4 U_g29816 ( .A1(g29759), .A2(g13883), .ZN(g29816) );
AND2_X4 U_g29817 ( .A1(g29709), .A2(g20694), .ZN(g29817) );
AND2_X4 U_g29818 ( .A1(g29732), .A2(g22293), .ZN(g29818) );
AND2_X4 U_g29819 ( .A1(g29751), .A2(g22294), .ZN(g29819) );
AND2_X4 U_g29820 ( .A1(g29717), .A2(g20743), .ZN(g29820) );
AND2_X4 U_g29821 ( .A1(g29731), .A2(g20746), .ZN(g29821) );
AND2_X4 U_g29822 ( .A1(g29705), .A2(g22335), .ZN(g29822) );
AND2_X4 U_g29827 ( .A1(g29741), .A2(g22356), .ZN(g29827) );
AND2_X4 U_g29828 ( .A1(g29740), .A2(g20802), .ZN(g29828) );
AND2_X4 U_g29833 ( .A1(g29725), .A2(g20813), .ZN(g29833) );
AND2_X4 U_g29834 ( .A1(g29713), .A2(g22366), .ZN(g29834) );
AND2_X4 U_g29839 ( .A1(g29747), .A2(g20827), .ZN(g29839) );
AND3_X4 U_g29909 ( .A1(g29735), .A2(g19420), .A3(g19401), .ZN(g29909) );
AND2_X4 U_g29910 ( .A1(g29779), .A2(g9961), .ZN(g29910) );
AND2_X4 U_g29942 ( .A1(g29771), .A2(g28877), .ZN(g29942) );
AND2_X4 U_g29944 ( .A1(g29782), .A2(g28889), .ZN(g29944) );
AND2_X4 U_g29945 ( .A1(g29773), .A2(g28894), .ZN(g29945) );
AND2_X4 U_g29946 ( .A1(g29778), .A2(g28906), .ZN(g29946) );
AND2_X4 U_g29947 ( .A1(g29785), .A2(g28911), .ZN(g29947) );
AND2_X4 U_g29948 ( .A1(g29775), .A2(g28916), .ZN(g29948) );
AND2_X4 U_g29949 ( .A1(g29781), .A2(g28932), .ZN(g29949) );
AND2_X4 U_g29950 ( .A1(g29788), .A2(g28937), .ZN(g29950) );
AND2_X4 U_g29951 ( .A1(g29777), .A2(g28945), .ZN(g29951) );
AND2_X4 U_g29952 ( .A1(g29784), .A2(g28959), .ZN(g29952) );
AND2_X4 U_g29953 ( .A1(g29791), .A2(g28967), .ZN(g29953) );
AND2_X4 U_g29954 ( .A1(g29770), .A2(g28975), .ZN(g29954) );
AND2_X4 U_g29955 ( .A1(g29787), .A2(g28993), .ZN(g29955) );
AND2_X4 U_g29956 ( .A1(g29780), .A2(g28998), .ZN(g29956) );
AND2_X4 U_g29957 ( .A1(g29772), .A2(g29005), .ZN(g29957) );
AND2_X4 U_g29958 ( .A1(g29783), .A2(g29027), .ZN(g29958) );
AND2_X4 U_g29959 ( .A1(g29774), .A2(g29035), .ZN(g29959) );
AND2_X4 U_g29960 ( .A1(g29786), .A2(g29050), .ZN(g29960) );
AND2_X4 U_g29961 ( .A1(g29776), .A2(g29057), .ZN(g29961) );
AND2_X4 U_g29962 ( .A1(g29789), .A2(g29069), .ZN(g29962) );
AND2_X4 U_g29963 ( .A1(g29758), .A2(g13737), .ZN(g29963) );
AND2_X4 U_g29964 ( .A1(g29757), .A2(g13786), .ZN(g29964) );
AND2_X4 U_g29965 ( .A1(g29756), .A2(g11961), .ZN(g29965) );
AND2_X4 U_g29966 ( .A1(g29755), .A2(g12004), .ZN(g29966) );
AND2_X4 U_g29967 ( .A1(g29754), .A2(g12066), .ZN(g29967) );
AND2_X4 U_g29968 ( .A1(g29765), .A2(g12119), .ZN(g29968) );
AND2_X4 U_g29969 ( .A1(g29721), .A2(g22237), .ZN(g29969) );
AND2_X4 U_g29970 ( .A1(g29764), .A2(g12178), .ZN(g29970) );
AND2_X4 U_g29971 ( .A1(g29763), .A2(g13861), .ZN(g29971) );
AND2_X4 U_g29980 ( .A1(g29881), .A2(g8324), .ZN(g29980) );
AND2_X4 U_g29981 ( .A1(g29869), .A2(g8330), .ZN(g29981) );
AND2_X4 U_g29982 ( .A1(g29893), .A2(g8336), .ZN(g29982) );
AND2_X4 U_g29983 ( .A1(g29885), .A2(g8344), .ZN(g29983) );
AND2_X4 U_g29984 ( .A1(g29873), .A2(g8351), .ZN(g29984) );
AND2_X4 U_g29985 ( .A1(g29897), .A2(g8363), .ZN(g29985) );
AND2_X4 U_g29986 ( .A1(g29877), .A2(g8366), .ZN(g29986) );
AND2_X4 U_g29987 ( .A1(g29889), .A2(g8369), .ZN(g29987) );
AND2_X4 U_g29988 ( .A1(g29881), .A2(g8382), .ZN(g29988) );
AND2_X4 U_g29989 ( .A1(g29893), .A2(g8391), .ZN(g29989) );
AND2_X4 U_g29990 ( .A1(g29885), .A2(g8397), .ZN(g29990) );
AND2_X4 U_g29991 ( .A1(g29901), .A2(g8403), .ZN(g29991) );
AND2_X4 U_g29992 ( .A1(g12441), .A2(g29909), .ZN(g29992) );
AND2_X4 U_g29993 ( .A1(g29897), .A2(g8411), .ZN(g29993) );
AND2_X4 U_g29994 ( .A1(g29889), .A2(g8418), .ZN(g29994) );
AND2_X4 U_g29995 ( .A1(g29893), .A2(g8434), .ZN(g29995) );
AND2_X4 U_g29996 ( .A1(g29901), .A2(g8443), .ZN(g29996) );
AND2_X4 U_g29997 ( .A1(g29918), .A2(g22277), .ZN(g29997) );
AND2_X4 U_g29998 ( .A1(g29922), .A2(g22278), .ZN(g29998) );
AND2_X4 U_g29999 ( .A1(g29924), .A2(g22279), .ZN(g29999) );
AND2_X4 U_g30000 ( .A1(g10767), .A2(g29930), .ZN(g30000) );
AND2_X4 U_g30001 ( .A1(g29897), .A2(g8449), .ZN(g30001) );
AND2_X4 U_g30002 ( .A1(g29905), .A2(g8455), .ZN(g30002) );
AND2_X4 U_g30003 ( .A1(g29901), .A2(g8469), .ZN(g30003) );
AND2_X4 U_g30004 ( .A1(g29926), .A2(g22295), .ZN(g30004) );
AND2_X4 U_g30005 ( .A1(g29905), .A2(g8478), .ZN(g30005) );
AND2_X4 U_g30006 ( .A1(g29928), .A2(g22310), .ZN(g30006) );
AND2_X4 U_g30007 ( .A1(g29905), .A2(g8494), .ZN(g30007) );
AND2_X4 U_g30008 ( .A1(g29919), .A2(g22334), .ZN(g30008) );
AND2_X4 U_g30009 ( .A1(g29929), .A2(g22357), .ZN(g30009) );
AND2_X4 U_g30077 ( .A1(g29823), .A2(g10963), .ZN(g30077) );
AND2_X4 U_g30079 ( .A1(g29823), .A2(g10988), .ZN(g30079) );
AND2_X4 U_g30080 ( .A1(g29829), .A2(g10996), .ZN(g30080) );
AND2_X4 U_g30081 ( .A1(g29823), .A2(g11022), .ZN(g30081) );
AND2_X4 U_g30082 ( .A1(g29829), .A2(g11036), .ZN(g30082) );
AND2_X4 U_g30083 ( .A1(g29835), .A2(g11048), .ZN(g30083) );
AND2_X4 U_g30085 ( .A1(g29829), .A2(g11092), .ZN(g30085) );
AND2_X4 U_g30086 ( .A1(g29835), .A2(g11108), .ZN(g30086) );
AND2_X4 U_g30087 ( .A1(g29840), .A2(g11120), .ZN(g30087) );
AND2_X4 U_g30088 ( .A1(g29844), .A2(g11138), .ZN(g30088) );
AND2_X4 U_g30089 ( .A1(g29835), .A2(g11160), .ZN(g30089) );
AND2_X4 U_g30090 ( .A1(g29840), .A2(g11176), .ZN(g30090) );
AND2_X4 U_g30091 ( .A1(g29844), .A2(g11202), .ZN(g30091) );
AND2_X4 U_g30092 ( .A1(g29849), .A2(g11205), .ZN(g30092) );
AND2_X4 U_g30093 ( .A1(g29853), .A2(g11222), .ZN(g30093) );
AND2_X4 U_g30094 ( .A1(g29840), .A2(g11246), .ZN(g30094) );
AND2_X4 U_g30095 ( .A1(g29857), .A2(g11265), .ZN(g30095) );
AND2_X4 U_g30096 ( .A1(g29844), .A2(g11268), .ZN(g30096) );
AND2_X4 U_g30097 ( .A1(g29849), .A2(g11271), .ZN(g30097) );
AND2_X4 U_g30098 ( .A1(g29853), .A2(g11284), .ZN(g30098) );
AND2_X4 U_g30099 ( .A1(g29861), .A2(g11287), .ZN(g30099) );
AND2_X4 U_g30100 ( .A1(g29865), .A2(g11306), .ZN(g30100) );
AND2_X4 U_g30101 ( .A1(g29857), .A2(g11341), .ZN(g30101) );
AND2_X4 U_g30102 ( .A1(g29849), .A2(g11348), .ZN(g30102) );
AND2_X4 U_g30103 ( .A1(g29869), .A2(g11358), .ZN(g30103) );
AND2_X4 U_g30104 ( .A1(g29853), .A2(g11361), .ZN(g30104) );
AND2_X4 U_g30105 ( .A1(g29861), .A2(g11364), .ZN(g30105) );
AND2_X4 U_g30106 ( .A1(g29865), .A2(g11379), .ZN(g30106) );
AND2_X4 U_g30107 ( .A1(g29873), .A2(g11382), .ZN(g30107) );
AND2_X4 U_g30108 ( .A1(g29877), .A2(g11401), .ZN(g30108) );
AND2_X4 U_g30109 ( .A1(g29857), .A2(g11411), .ZN(g30109) );
AND2_X4 U_g30110 ( .A1(g29881), .A2(g11417), .ZN(g30110) );
AND2_X4 U_g30111 ( .A1(g29869), .A2(g11425), .ZN(g30111) );
AND2_X4 U_g30112 ( .A1(g29861), .A2(g11432), .ZN(g30112) );
AND2_X4 U_g30113 ( .A1(g29885), .A2(g11444), .ZN(g30113) );
AND2_X4 U_g30114 ( .A1(g29865), .A2(g11447), .ZN(g30114) );
AND2_X4 U_g30115 ( .A1(g29873), .A2(g11450), .ZN(g30115) );
AND2_X4 U_g30116 ( .A1(g29921), .A2(g22236), .ZN(g30116) );
AND2_X4 U_g30117 ( .A1(g29877), .A2(g11465), .ZN(g30117) );
AND2_X4 U_g30118 ( .A1(g29889), .A2(g11468), .ZN(g30118) );
AND2_X4 U_g30123 ( .A1(g30070), .A2(g20641), .ZN(g30123) );
AND2_X4 U_g30127 ( .A1(g30065), .A2(g20719), .ZN(g30127) );
AND2_X4 U_g30128 ( .A1(g30062), .A2(g20722), .ZN(g30128) );
AND2_X4 U_g30129 ( .A1(g30071), .A2(g20725), .ZN(g30129) );
AND2_X4 U_g30131 ( .A1(g30059), .A2(g20749), .ZN(g30131) );
AND2_X4 U_g30132 ( .A1(g30068), .A2(g20776), .ZN(g30132) );
AND2_X4 U_g30133 ( .A1(g30067), .A2(g20799), .ZN(g30133) );
AND2_X4 U_g30138 ( .A1(g30069), .A2(g20816), .ZN(g30138) );
AND2_X4 U_g30216 ( .A1(g30036), .A2(g8921), .ZN(g30216) );
AND2_X4 U_g30217 ( .A1(g30036), .A2(g8955), .ZN(g30217) );
AND2_X4 U_g30218 ( .A1(g30040), .A2(g8961), .ZN(g30218) );
AND2_X4 U_g30219 ( .A1(g30036), .A2(g8980), .ZN(g30219) );
AND2_X4 U_g30220 ( .A1(g30040), .A2(g8987), .ZN(g30220) );
AND2_X4 U_g30221 ( .A1(g30044), .A2(g8993), .ZN(g30221) );
AND2_X4 U_g30222 ( .A1(g30040), .A2(g9010), .ZN(g30222) );
AND2_X4 U_g30223 ( .A1(g30044), .A2(g9016), .ZN(g30223) );
AND2_X4 U_g30224 ( .A1(g30048), .A2(g9022), .ZN(g30224) );
AND2_X4 U_g30225 ( .A1(g30044), .A2(g9035), .ZN(g30225) );
AND2_X4 U_g30226 ( .A1(g30048), .A2(g9041), .ZN(g30226) );
AND2_X4 U_g30227 ( .A1(g30048), .A2(g9058), .ZN(g30227) );
AND2_X4 U_g30327 ( .A1(g30187), .A2(g8321), .ZN(g30327) );
AND2_X4 U_g30330 ( .A1(g30195), .A2(g8333), .ZN(g30330) );
AND2_X4 U_g30333 ( .A1(g30191), .A2(g8341), .ZN(g30333) );
AND2_X4 U_g30334 ( .A1(g30203), .A2(g8347), .ZN(g30334) );
AND2_X4 U_g30337 ( .A1(g30199), .A2(g8354), .ZN(g30337) );
AND2_X4 U_g30340 ( .A1(g30207), .A2(g8372), .ZN(g30340) );
AND2_X4 U_g30345 ( .A1(g30195), .A2(g8388), .ZN(g30345) );
AND2_X4 U_g30348 ( .A1(g30203), .A2(g8400), .ZN(g30348) );
AND2_X4 U_g30351 ( .A1(g30199), .A2(g8408), .ZN(g30351) );
AND2_X4 U_g30352 ( .A1(g30211), .A2(g8414), .ZN(g30352) );
AND2_X4 U_g30355 ( .A1(g30207), .A2(g8421), .ZN(g30355) );
AND2_X4 U_g30361 ( .A1(g30203), .A2(g8440), .ZN(g30361) );
AND2_X4 U_g30364 ( .A1(g30211), .A2(g8452), .ZN(g30364) );
AND2_X4 U_g30367 ( .A1(g30207), .A2(g8460), .ZN(g30367) );
AND2_X4 U_g30372 ( .A1(g8594), .A2(g30228), .ZN(g30372) );
AND2_X4 U_g30374 ( .A1(g30211), .A2(g8475), .ZN(g30374) );
AND2_X4 U_g30387 ( .A1(g30229), .A2(g8888), .ZN(g30387) );
AND2_X4 U_g30388 ( .A1(g30229), .A2(g8918), .ZN(g30388) );
AND2_X4 U_g30389 ( .A1(g30233), .A2(g8928), .ZN(g30389) );
AND2_X4 U_g30390 ( .A1(g30229), .A2(g8952), .ZN(g30390) );
AND2_X4 U_g30391 ( .A1(g30233), .A2(g8958), .ZN(g30391) );
AND2_X4 U_g30392 ( .A1(g30237), .A2(g8968), .ZN(g30392) );
AND2_X4 U_g30393 ( .A1(g30233), .A2(g8984), .ZN(g30393) );
AND2_X4 U_g30394 ( .A1(g30237), .A2(g8990), .ZN(g30394) );
AND2_X4 U_g30395 ( .A1(g30241), .A2(g9000), .ZN(g30395) );
AND2_X4 U_g30396 ( .A1(g30237), .A2(g9013), .ZN(g30396) );
AND2_X4 U_g30397 ( .A1(g30241), .A2(g9019), .ZN(g30397) );
AND2_X4 U_g30398 ( .A1(g30241), .A2(g9038), .ZN(g30398) );
AND2_X4 U_g30407 ( .A1(g30134), .A2(g10991), .ZN(g30407) );
AND2_X4 U_g30409 ( .A1(g30134), .A2(g11025), .ZN(g30409) );
AND2_X4 U_g30410 ( .A1(g30139), .A2(g11028), .ZN(g30410) );
AND2_X4 U_g30411 ( .A1(g30143), .A2(g11039), .ZN(g30411) );
AND2_X4 U_g30436 ( .A1(g30134), .A2(g11079), .ZN(g30436) );
AND2_X4 U_g30437 ( .A1(g30139), .A2(g11082), .ZN(g30437) );
AND2_X4 U_g30438 ( .A1(g30147), .A2(g11085), .ZN(g30438) );
AND2_X4 U_g30440 ( .A1(g30143), .A2(g11095), .ZN(g30440) );
AND2_X4 U_g30441 ( .A1(g30151), .A2(g11098), .ZN(g30441) );
AND2_X4 U_g30442 ( .A1(g30155), .A2(g11111), .ZN(g30442) );
AND2_X4 U_g30444 ( .A1(g30139), .A2(g11132), .ZN(g30444) );
AND2_X4 U_g30445 ( .A1(g30147), .A2(g11135), .ZN(g30445) );
AND2_X4 U_g30447 ( .A1(g30143), .A2(g11145), .ZN(g30447) );
AND2_X4 U_g30448 ( .A1(g30151), .A2(g11148), .ZN(g30448) );
AND2_X4 U_g30449 ( .A1(g30159), .A2(g11151), .ZN(g30449) );
AND2_X4 U_g30451 ( .A1(g30155), .A2(g11163), .ZN(g30451) );
AND2_X4 U_g30452 ( .A1(g30163), .A2(g11166), .ZN(g30452) );
AND2_X4 U_g30453 ( .A1(g30167), .A2(g11179), .ZN(g30453) );
AND2_X4 U_g30454 ( .A1(g30147), .A2(g11199), .ZN(g30454) );
AND2_X4 U_g30457 ( .A1(g30151), .A2(g11216), .ZN(g30457) );
AND2_X4 U_g30458 ( .A1(g30159), .A2(g11219), .ZN(g30458) );
AND2_X4 U_g30460 ( .A1(g30155), .A2(g11231), .ZN(g30460) );
AND2_X4 U_g30461 ( .A1(g30163), .A2(g11234), .ZN(g30461) );
AND2_X4 U_g30462 ( .A1(g30171), .A2(g11237), .ZN(g30462) );
AND2_X4 U_g30464 ( .A1(g30167), .A2(g11249), .ZN(g30464) );
AND2_X4 U_g30465 ( .A1(g30175), .A2(g11252), .ZN(g30465) );
AND2_X4 U_g30467 ( .A1(g30179), .A2(g11274), .ZN(g30467) );
AND2_X4 U_g30469 ( .A1(g30159), .A2(g11281), .ZN(g30469) );
AND2_X4 U_g30472 ( .A1(g30163), .A2(g11300), .ZN(g30472) );
AND2_X4 U_g30473 ( .A1(g30171), .A2(g11303), .ZN(g30473) );
AND2_X4 U_g30475 ( .A1(g30167), .A2(g11315), .ZN(g30475) );
AND2_X4 U_g30476 ( .A1(g30175), .A2(g11318), .ZN(g30476) );
AND2_X4 U_g30477 ( .A1(g30183), .A2(g11321), .ZN(g30477) );
AND2_X4 U_g30478 ( .A1(g30187), .A2(g11344), .ZN(g30478) );
AND2_X4 U_g30481 ( .A1(g30179), .A2(g11351), .ZN(g30481) );
AND2_X4 U_g30484 ( .A1(g30191), .A2(g11367), .ZN(g30484) );
AND2_X4 U_g30486 ( .A1(g30171), .A2(g11376), .ZN(g30486) );
AND2_X4 U_g30489 ( .A1(g30175), .A2(g11395), .ZN(g30489) );
AND2_X4 U_g30490 ( .A1(g30183), .A2(g11398), .ZN(g30490) );
AND2_X4 U_g30492 ( .A1(g30187), .A2(g11414), .ZN(g30492) );
AND2_X4 U_g30495 ( .A1(g30179), .A2(g11422), .ZN(g30495) );
AND2_X4 U_g30496 ( .A1(g30195), .A2(g11428), .ZN(g30496) );
AND2_X4 U_g30499 ( .A1(g30191), .A2(g11435), .ZN(g30499) );
AND2_X4 U_g30502 ( .A1(g30199), .A2(g11453), .ZN(g30502) );
AND2_X4 U_g30504 ( .A1(g30183), .A2(g11462), .ZN(g30504) );
AND2_X4 U_g30696 ( .A1(g30383), .A2(g10943), .ZN(g30696) );
AND2_X4 U_g30697 ( .A1(g30383), .A2(g11011), .ZN(g30697) );
AND2_X4 U_g30698 ( .A1(g30383), .A2(g11126), .ZN(g30698) );
AND2_X4 U_g30728 ( .A1(g30605), .A2(g22252), .ZN(g30728) );
AND2_X4 U_g30735 ( .A1(g30629), .A2(g22268), .ZN(g30735) );
AND2_X4 U_g30736 ( .A1(g30584), .A2(g20669), .ZN(g30736) );
AND2_X4 U_g30743 ( .A1(g30610), .A2(g22283), .ZN(g30743) );
AND2_X4 U_g30744 ( .A1(g30609), .A2(g20697), .ZN(g30744) );
AND2_X4 U_g30750 ( .A1(g30593), .A2(g20729), .ZN(g30750) );
AND2_X4 U_g30754 ( .A1(g30614), .A2(g22313), .ZN(g30754) );
AND2_X4 U_g30755 ( .A1(g30632), .A2(g22314), .ZN(g30755) );
AND2_X4 U_g30757 ( .A1(g30601), .A2(g20780), .ZN(g30757) );
AND2_X4 U_g30758 ( .A1(g30613), .A2(g20783), .ZN(g30758) );
AND2_X4 U_g30759 ( .A1(g30588), .A2(g22360), .ZN(g30759) );
AND2_X4 U_g30760 ( .A1(g30622), .A2(g22379), .ZN(g30760) );
AND2_X4 U_g30761 ( .A1(g30621), .A2(g20822), .ZN(g30761) );
AND2_X4 U_g30762 ( .A1(g30608), .A2(g20830), .ZN(g30762) );
AND2_X4 U_g30763 ( .A1(g30597), .A2(g22386), .ZN(g30763) );
AND2_X4 U_g30764 ( .A1(g30628), .A2(g20837), .ZN(g30764) );
AND3_X4 U_g30766 ( .A1(g30617), .A2(g19457), .A3(g19431), .ZN(g30766) );
AND2_X4 U_g30916 ( .A1(g30785), .A2(g22251), .ZN(g30916) );
AND2_X4 U_g30917 ( .A1(g12446), .A2(g30766), .ZN(g30917) );
AND2_X4 U_g30918 ( .A1(g30780), .A2(g22296), .ZN(g30918) );
AND2_X4 U_g30919 ( .A1(g30786), .A2(g22297), .ZN(g30919) );
AND2_X4 U_g30920 ( .A1(g30787), .A2(g22298), .ZN(g30920) );
AND2_X4 U_g30921 ( .A1(g10773), .A2(g30791), .ZN(g30921) );
AND2_X4 U_g30922 ( .A1(g30788), .A2(g22315), .ZN(g30922) );
AND2_X4 U_g30923 ( .A1(g30789), .A2(g22338), .ZN(g30923) );
AND2_X4 U_g30924 ( .A1(g30783), .A2(g22359), .ZN(g30924) );
AND2_X4 U_g30925 ( .A1(g30790), .A2(g22380), .ZN(g30925) );
AND2_X4 U_g30944 ( .A1(g30935), .A2(g20666), .ZN(g30944) );
AND2_X4 U_g30945 ( .A1(g30931), .A2(g20754), .ZN(g30945) );
AND2_X4 U_g30946 ( .A1(g30930), .A2(g20757), .ZN(g30946) );
AND2_X4 U_g30947 ( .A1(g30936), .A2(g20760), .ZN(g30947) );
AND2_X4 U_g30948 ( .A1(g30929), .A2(g20786), .ZN(g30948) );
AND2_X4 U_g30949 ( .A1(g30933), .A2(g20806), .ZN(g30949) );
AND2_X4 U_g30950 ( .A1(g30932), .A2(g20819), .ZN(g30950) );
AND2_X4 U_g30951 ( .A1(g30934), .A2(g20833), .ZN(g30951) );
AND2_X4 U_g30953 ( .A1(g8605), .A2(g30952), .ZN(g30953) );
OR2_X4 U_g9144 ( .A1(g2986), .A2(g5389), .ZN(g9144) );
OR2_X4 U_g10778 ( .A1(g2929), .A2(g8022), .ZN(g10778) );
OR2_X4 U_g12377 ( .A1(g7553), .A2(g11059), .ZN(g12377) );
OR2_X4 U_g12407 ( .A1(g7573), .A2(g10779), .ZN(g12407) );
OR2_X4 U_g12886 ( .A1(g9534), .A2(g3398), .ZN(g12886) );
OR2_X4 U_g12926 ( .A1(g9676), .A2(g3554), .ZN(g12926) );
OR2_X4 U_g12955 ( .A1(g9822), .A2(g3710), .ZN(g12955) );
OR2_X4 U_g12984 ( .A1(g9968), .A2(g3866), .ZN(g12984) );
OR2_X4 U_g16539 ( .A1(g15880), .A2(g14657), .ZN(g16539) );
OR2_X4 U_g16571 ( .A1(g15913), .A2(g14691), .ZN(g16571) );
OR2_X4 U_g16595 ( .A1(g15942), .A2(g14725), .ZN(g16595) );
OR2_X4 U_g16615 ( .A1(g15971), .A2(g14753), .ZN(g16615) );
OR2_X4 U_g17973 ( .A1(g11623), .A2(g15659), .ZN(g17973) );
OR2_X4 U_g19181 ( .A1(g17729), .A2(g17979), .ZN(g19181) );
OR2_X4 U_g19186 ( .A1(g18419), .A2(g17887), .ZN(g19186) );
OR2_X4 U_g19187 ( .A1(g18419), .A2(g17729), .ZN(g19187) );
OR2_X4 U_g19188 ( .A1(g17830), .A2(g18096), .ZN(g19188) );
OR2_X4 U_g19191 ( .A1(g17807), .A2(g17887), .ZN(g19191) );
OR2_X4 U_g19192 ( .A1(g18183), .A2(g18270), .ZN(g19192) );
OR2_X4 U_g19193 ( .A1(g18492), .A2(g17998), .ZN(g19193) );
OR2_X4 U_g19194 ( .A1(g18492), .A2(g17830), .ZN(g19194) );
OR2_X4 U_g19195 ( .A1(g17942), .A2(g18212), .ZN(g19195) );
OR2_X4 U_g19200 ( .A1(g18346), .A2(g18424), .ZN(g19200) );
OR2_X4 U_g19201 ( .A1(g18183), .A2(g18424), .ZN(g19201) );
OR2_X4 U_g19202 ( .A1(g17919), .A2(g17998), .ZN(g19202) );
OR2_X4 U_g19203 ( .A1(g18290), .A2(g18363), .ZN(g19203) );
OR2_X4 U_g19204 ( .A1(g18556), .A2(g18115), .ZN(g19204) );
OR2_X4 U_g19205 ( .A1(g18556), .A2(g17942), .ZN(g19205) );
OR2_X4 U_g19206 ( .A1(g18053), .A2(g18319), .ZN(g19206) );
OR2_X4 U_g19209 ( .A1(g18079), .A2(g18346), .ZN(g19209) );
OR2_X4 U_g19210 ( .A1(g18079), .A2(g18183), .ZN(g19210) );
OR2_X4 U_g19211 ( .A1(g18441), .A2(g18497), .ZN(g19211) );
OR2_X4 U_g19212 ( .A1(g18290), .A2(g18497), .ZN(g19212) );
OR2_X4 U_g19213 ( .A1(g18030), .A2(g18115), .ZN(g19213) );
OR2_X4 U_g19214 ( .A1(g18383), .A2(g18458), .ZN(g19214) );
OR2_X4 U_g19215 ( .A1(g18606), .A2(g18231), .ZN(g19215) );
OR2_X4 U_g19216 ( .A1(g18606), .A2(g18053), .ZN(g19216) );
OR2_X4 U_g19221 ( .A1(g18270), .A2(g18346), .ZN(g19221) );
OR2_X4 U_g19222 ( .A1(g18195), .A2(g18441), .ZN(g19222) );
OR2_X4 U_g19223 ( .A1(g18195), .A2(g18290), .ZN(g19223) );
OR2_X4 U_g19224 ( .A1(g18514), .A2(g18561), .ZN(g19224) );
OR2_X4 U_g19225 ( .A1(g18383), .A2(g18561), .ZN(g19225) );
OR2_X4 U_g19226 ( .A1(g18147), .A2(g18231), .ZN(g19226) );
OR2_X4 U_g19227 ( .A1(g18478), .A2(g18531), .ZN(g19227) );
OR3_X4 U_I25477 ( .A1(g17024), .A2(g17000), .A3(g16992), .ZN(I25477) );
OR3_X4 U_g19230 ( .A1(g16985), .A2(g16965), .A3(I25477), .ZN(g19230) );
OR2_X4 U_g19231 ( .A1(g18363), .A2(g18441), .ZN(g19231) );
OR2_X4 U_g19232 ( .A1(g18302), .A2(g18514), .ZN(g19232) );
OR2_X4 U_g19233 ( .A1(g18302), .A2(g18383), .ZN(g19233) );
OR2_X4 U_g19234 ( .A1(g18578), .A2(g18611), .ZN(g19234) );
OR2_X4 U_g19235 ( .A1(g18478), .A2(g18611), .ZN(g19235) );
OR3_X4 U_I25495 ( .A1(g17158), .A2(g17137), .A3(g17115), .ZN(I25495) );
OR3_X4 U_g19240 ( .A1(g17083), .A2(g17050), .A3(I25495), .ZN(g19240) );
OR2_X4 U_g19242 ( .A1(g14244), .A2(g16501), .ZN(g19242) );
OR3_X4 U_I25500 ( .A1(g17058), .A2(g17030), .A3(g17016), .ZN(I25500) );
OR3_X4 U_g19243 ( .A1(g16995), .A2(g16986), .A3(I25500), .ZN(g19243) );
OR2_X4 U_g19244 ( .A1(g18458), .A2(g18514), .ZN(g19244) );
OR2_X4 U_g19245 ( .A1(g18395), .A2(g18578), .ZN(g19245) );
OR2_X4 U_g19246 ( .A1(g18395), .A2(g18478), .ZN(g19246) );
OR2_X4 U_g19250 ( .A1(g17729), .A2(g17807), .ZN(g19250) );
OR3_X4 U_I25516 ( .A1(g17173), .A2(g17160), .A3(g17142), .ZN(I25516) );
OR3_X4 U_g19253 ( .A1(g17121), .A2(g17085), .A3(I25516), .ZN(g19253) );
OR2_X4 U_g19255 ( .A1(g14366), .A2(g16523), .ZN(g19255) );
OR3_X4 U_I25521 ( .A1(g17093), .A2(g17064), .A3(g17046), .ZN(I25521) );
OR3_X4 U_g19256 ( .A1(g17019), .A2(g16996), .A3(I25521), .ZN(g19256) );
OR2_X4 U_g19257 ( .A1(g18531), .A2(g18578), .ZN(g19257) );
OR2_X4 U_g19263 ( .A1(g17887), .A2(g17979), .ZN(g19263) );
OR2_X4 U_g19264 ( .A1(g17830), .A2(g17919), .ZN(g19264) );
OR3_X4 U_I25549 ( .A1(g17190), .A2(g17175), .A3(g17165), .ZN(I25549) );
OR3_X4 U_g19266 ( .A1(g17148), .A2(g17123), .A3(I25549), .ZN(g19266) );
OR2_X4 U_g19268 ( .A1(g14478), .A2(g16554), .ZN(g19268) );
OR3_X4 U_I25554 ( .A1(g17131), .A2(g17099), .A3(g17080), .ZN(I25554) );
OR3_X4 U_g19269 ( .A1(g17049), .A2(g17020), .A3(I25554), .ZN(g19269) );
OR3_X4 U_g19275 ( .A1(g16867), .A2(g16515), .A3(g19001), .ZN(g19275) );
OR2_X4 U_g19278 ( .A1(g17998), .A2(g18096), .ZN(g19278) );
OR2_X4 U_g19279 ( .A1(g17942), .A2(g18030), .ZN(g19279) );
OR3_X4 U_I25588 ( .A1(g17201), .A2(g17192), .A3(g17180), .ZN(I25588) );
OR3_X4 U_g19281 ( .A1(g17171), .A2(g17150), .A3(I25588), .ZN(g19281) );
OR2_X4 U_g19283 ( .A1(g14565), .A2(g16586), .ZN(g19283) );
OR3_X4 U_g19294 ( .A1(g16895), .A2(g16546), .A3(g16507), .ZN(g19294) );
OR2_X4 U_g19297 ( .A1(g18115), .A2(g18212), .ZN(g19297) );
OR2_X4 U_g19298 ( .A1(g18053), .A2(g18147), .ZN(g19298) );
OR3_X4 U_g19312 ( .A1(g16924), .A2(g16578), .A3(g16529), .ZN(g19312) );
OR2_X4 U_g19315 ( .A1(g18231), .A2(g18319), .ZN(g19315) );
OR3_X4 U_g19333 ( .A1(g16954), .A2(g16602), .A3(g16560), .ZN(g19333) );
OR2_X4 U_g19450 ( .A1(g14837), .A2(g16682), .ZN(g19450) );
OR2_X4 U_g19477 ( .A1(g14910), .A2(g16708), .ZN(g19477) );
OR2_X4 U_g19500 ( .A1(g14991), .A2(g16739), .ZN(g19500) );
OR3_X4 U_g19503 ( .A1(g16884), .A2(g16697), .A3(g16665), .ZN(g19503) );
OR2_X4 U_g19521 ( .A1(g15080), .A2(g16781), .ZN(g19521) );
OR3_X4 U_g19522 ( .A1(g16913), .A2(g16728), .A3(g16686), .ZN(g19522) );
OR3_X4 U_g19532 ( .A1(g16943), .A2(g16770), .A3(g16712), .ZN(g19532) );
OR3_X4 U_g19542 ( .A1(g16974), .A2(g16797), .A3(g16743), .ZN(g19542) );
OR3_X4 U_I26429 ( .A1(g17979), .A2(g17887), .A3(g17807), .ZN(I26429) );
OR3_X4 U_g19981 ( .A1(g17729), .A2(g18419), .A3(I26429), .ZN(g19981) );
OR3_X4 U_I26455 ( .A1(g18424), .A2(g18346), .A3(g18270), .ZN(I26455) );
OR3_X4 U_g20015 ( .A1(g18183), .A2(g18079), .A3(I26455), .ZN(g20015) );
OR3_X4 U_I26461 ( .A1(g18096), .A2(g17998), .A3(g17919), .ZN(I26461) );
OR3_X4 U_g20019 ( .A1(g17830), .A2(g18492), .A3(I26461), .ZN(g20019) );
OR3_X4 U_I26491 ( .A1(g18497), .A2(g18441), .A3(g18363), .ZN(I26491) );
OR3_X4 U_g20057 ( .A1(g18290), .A2(g18195), .A3(I26491), .ZN(g20057) );
OR3_X4 U_I26497 ( .A1(g18212), .A2(g18115), .A3(g18030), .ZN(I26497) );
OR3_X4 U_g20061 ( .A1(g17942), .A2(g18556), .A3(I26497), .ZN(g20061) );
OR3_X4 U_I26532 ( .A1(g18561), .A2(g18514), .A3(g18458), .ZN(I26532) );
OR3_X4 U_g20098 ( .A1(g18383), .A2(g18302), .A3(I26532), .ZN(g20098) );
OR3_X4 U_I26538 ( .A1(g18319), .A2(g18231), .A3(g18147), .ZN(I26538) );
OR3_X4 U_g20102 ( .A1(g18053), .A2(g18606), .A3(I26538), .ZN(g20102) );
OR3_X4 U_I26571 ( .A1(g18611), .A2(g18578), .A3(g18531), .ZN(I26571) );
OR3_X4 U_g20123 ( .A1(g18478), .A2(g18395), .A3(I26571), .ZN(g20123) );
OR3_X4 U_g21120 ( .A1(g19484), .A2(g16515), .A3(g14071), .ZN(g21120) );
OR3_X4 U_g21139 ( .A1(g19505), .A2(g16546), .A3(g14186), .ZN(g21139) );
OR3_X4 U_g21159 ( .A1(g19524), .A2(g16578), .A3(g14301), .ZN(g21159) );
OR3_X4 U_g21179 ( .A1(g19534), .A2(g16602), .A3(g14423), .ZN(g21179) );
OR3_X4 U_g21244 ( .A1(g19578), .A2(g16697), .A3(g14776), .ZN(g21244) );
OR3_X4 U_g21253 ( .A1(g19608), .A2(g16728), .A3(g14811), .ZN(g21253) );
OR3_X4 U_g21261 ( .A1(g19641), .A2(g16770), .A3(g14863), .ZN(g21261) );
OR3_X4 U_g21269 ( .A1(g19681), .A2(g16797), .A3(g14936), .ZN(g21269) );
OR3_X4 U_g21501 ( .A1(g20522), .A2(g16867), .A3(g14071), .ZN(g21501) );
OR3_X4 U_g21536 ( .A1(g20522), .A2(g19484), .A3(g19001), .ZN(g21536) );
OR3_X4 U_g21540 ( .A1(g20542), .A2(g16895), .A3(g14186), .ZN(g21540) );
OR3_X4 U_g21572 ( .A1(g20542), .A2(g19505), .A3(g16507), .ZN(g21572) );
OR3_X4 U_g21576 ( .A1(g19067), .A2(g16924), .A3(g14301), .ZN(g21576) );
OR3_X4 U_g21605 ( .A1(g19067), .A2(g19524), .A3(g16529), .ZN(g21605) );
OR3_X4 U_g21609 ( .A1(g19084), .A2(g16954), .A3(g14423), .ZN(g21609) );
OR3_X4 U_g21634 ( .A1(g19084), .A2(g19534), .A3(g16560), .ZN(g21634) );
OR3_X4 U_g21774 ( .A1(g19121), .A2(g16884), .A3(g14776), .ZN(g21774) );
OR3_X4 U_g21787 ( .A1(g19121), .A2(g19578), .A3(g16665), .ZN(g21787) );
OR3_X4 U_I28305 ( .A1(g20197), .A2(g20177), .A3(g20145), .ZN(I28305) );
OR3_X4 U_g21788 ( .A1(g20117), .A2(g20094), .A3(I28305), .ZN(g21788) );
OR3_X4 U_g21789 ( .A1(g19128), .A2(g16913), .A3(g14811), .ZN(g21789) );
OR3_X4 U_I28318 ( .A1(g19092), .A2(g19088), .A3(g19079), .ZN(I28318) );
OR4_X4 U_g21799 ( .A1(g16505), .A2(g20538), .A3(g18994), .A4(I28318), .ZN(g21799) );
OR4_X4 U_g21800 ( .A1(g18665), .A2(g20270), .A3(g20248), .A4(g18647), .ZN(g21800) );
OR3_X4 U_g21801 ( .A1(g19128), .A2(g19608), .A3(g16686), .ZN(g21801) );
OR3_X4 U_I28323 ( .A1(g20227), .A2(g20211), .A3(g20183), .ZN(I28323) );
OR3_X4 U_g21802 ( .A1(g20147), .A2(g20119), .A3(I28323), .ZN(g21802) );
OR3_X4 U_g21803 ( .A1(g19135), .A2(g16943), .A3(g14863), .ZN(g21803) );
OR4_X4 U_g21806 ( .A1(g20116), .A2(g20093), .A3(g18547), .A4(g19097), .ZN(g21806) );
OR3_X4 U_I28330 ( .A1(g19099), .A2(g19094), .A3(g19089), .ZN(I28330) );
OR4_X4 U_g21807 ( .A1(g16527), .A2(g19063), .A3(g19007), .A4(I28330), .ZN(g21807) );
OR4_X4 U_g21808 ( .A1(g18688), .A2(g20282), .A3(g20271), .A4(g18650), .ZN(g21808) );
OR3_X4 U_g21809 ( .A1(g19135), .A2(g19641), .A3(g16712), .ZN(g21809) );
OR3_X4 U_I28335 ( .A1(g20254), .A2(g20241), .A3(g20217), .ZN(I28335) );
OR3_X4 U_g21810 ( .A1(g20185), .A2(g20149), .A3(I28335), .ZN(g21810) );
OR3_X4 U_g21811 ( .A1(g19138), .A2(g16974), .A3(g14936), .ZN(g21811) );
OR4_X4 U_g21813 ( .A1(g20146), .A2(g20118), .A3(g18597), .A4(g19104), .ZN(g21813) );
OR3_X4 U_I28341 ( .A1(g19106), .A2(g19101), .A3(g19095), .ZN(I28341) );
OR4_X4 U_g21814 ( .A1(g16558), .A2(g19080), .A3(g16513), .A4(I28341), .ZN(g21814) );
OR4_X4 U_g21815 ( .A1(g18717), .A2(g20293), .A3(g20283), .A4(g18654), .ZN(g21815) );
OR3_X4 U_g21816 ( .A1(g19138), .A2(g19681), .A3(g16743), .ZN(g21816) );
OR3_X4 U_I28346 ( .A1(g20277), .A2(g20268), .A3(g20247), .ZN(I28346) );
OR3_X4 U_g21817 ( .A1(g20219), .A2(g20187), .A3(I28346), .ZN(g21817) );
OR4_X4 U_g21819 ( .A1(g20184), .A2(g20148), .A3(g18629), .A4(g19109), .ZN(g21819) );
OR3_X4 U_I28351 ( .A1(g19111), .A2(g19108), .A3(g19102), .ZN(I28351) );
OR4_X4 U_g21820 ( .A1(g16590), .A2(g19090), .A3(g16535), .A4(I28351), .ZN(g21820) );
OR4_X4 U_g21821 ( .A1(g18753), .A2(g20309), .A3(g20294), .A4(g18668), .ZN(g21821) );
OR4_X4 U_g21823 ( .A1(g20218), .A2(g20186), .A3(g18638), .A4(g19116), .ZN(g21823) );
OR3_X4 U_I28365 ( .A1(g20280), .A2(g18652), .A3(g18649), .ZN(I28365) );
OR3_X4 U_g21844 ( .A1(g20222), .A2(g18645), .A3(I28365), .ZN(g21844) );
OR3_X4 U_I28369 ( .A1(g20291), .A2(g18666), .A3(g18653), .ZN(I28369) );
OR3_X4 U_g21846 ( .A1(g20249), .A2(g18648), .A3(I28369), .ZN(g21846) );
OR3_X4 U_I28374 ( .A1(g20307), .A2(g18689), .A3(g18667), .ZN(I28374) );
OR3_X4 U_g21849 ( .A1(g20272), .A2(g18651), .A3(I28374), .ZN(g21849) );
OR3_X4 U_I28380 ( .A1(g20326), .A2(g18718), .A3(g18690), .ZN(I28380) );
OR3_X4 U_g21856 ( .A1(g20284), .A2(g18655), .A3(I28380), .ZN(g21856) );
OR2_X4 U_g22175 ( .A1(g16075), .A2(g20842), .ZN(g22175) );
OR2_X4 U_g22190 ( .A1(g16113), .A2(g20850), .ZN(g22190) );
OR2_X4 U_g22199 ( .A1(g16164), .A2(g20858), .ZN(g22199) );
OR2_X4 U_g22205 ( .A1(g16223), .A2(g20866), .ZN(g22205) );
OR4_X4 U_g22811 ( .A1(g562), .A2(g559), .A3(g12451), .A4(g21851), .ZN(g22811) );
OR3_X4 U_g23052 ( .A1(g21800), .A2(g21788), .A3(g21844), .ZN(g23052) );
OR3_X4 U_g23071 ( .A1(g21808), .A2(g21802), .A3(g21846), .ZN(g23071) );
OR3_X4 U_g23084 ( .A1(g21815), .A2(g21810), .A3(g21849), .ZN(g23084) );
OR2_X4 U_g23089 ( .A1(g21806), .A2(g21799), .ZN(g23089) );
OR3_X4 U_g23100 ( .A1(g21821), .A2(g21817), .A3(g21856), .ZN(g23100) );
OR2_X4 U_g23107 ( .A1(g21813), .A2(g21807), .ZN(g23107) );
OR2_X4 U_g23120 ( .A1(g21819), .A2(g21814), .ZN(g23120) );
OR2_X4 U_g23129 ( .A1(g21823), .A2(g21820), .ZN(g23129) );
OR2_X4 U_g23319 ( .A1(g14493), .A2(g22385), .ZN(g23319) );
OR2_X4 U_g23688 ( .A1(g23106), .A2(g21906), .ZN(g23688) );
OR2_X4 U_g23742 ( .A1(g23119), .A2(g21920), .ZN(g23742) );
OR2_X4 U_g23797 ( .A1(g23128), .A2(g21938), .ZN(g23797) );
OR2_X4 U_g23850 ( .A1(g23139), .A2(g20647), .ZN(g23850) );
OR2_X4 U_g23919 ( .A1(g22666), .A2(g23140), .ZN(g23919) );
OR2_X4 U_g24239 ( .A1(g19387), .A2(g22401), .ZN(g24239) );
OR2_X4 U_g24244 ( .A1(g14144), .A2(g22317), .ZN(g24244) );
OR2_X4 U_g24245 ( .A1(g19417), .A2(g22402), .ZN(g24245) );
OR2_X4 U_g24252 ( .A1(g14259), .A2(g22342), .ZN(g24252) );
OR2_X4 U_g24254 ( .A1(g19454), .A2(g22403), .ZN(g24254) );
OR2_X4 U_g24257 ( .A1(g14381), .A2(g22365), .ZN(g24257) );
OR2_X4 U_g24258 ( .A1(g19481), .A2(g22404), .ZN(g24258) );
OR2_X4 U_g24633 ( .A1(g24094), .A2(g20842), .ZN(g24633) );
OR2_X4 U_g24653 ( .A1(g24095), .A2(g20850), .ZN(g24653) );
OR2_X4 U_g24672 ( .A1(g24097), .A2(g20858), .ZN(g24672) );
OR2_X4 U_g24691 ( .A1(g24103), .A2(g20866), .ZN(g24691) );
OR2_X4 U_g24890 ( .A1(g23639), .A2(g23144), .ZN(g24890) );
OR2_X4 U_g24909 ( .A1(g23726), .A2(g23142), .ZN(g24909) );
OR2_X4 U_g24925 ( .A1(g23772), .A2(g23141), .ZN(g24925) );
OR2_X4 U_g24965 ( .A1(g23922), .A2(g23945), .ZN(g24965) );
OR2_X4 U_g24978 ( .A1(g23954), .A2(g23974), .ZN(g24978) );
OR2_X4 U_g24989 ( .A1(g23983), .A2(g24004), .ZN(g24989) );
OR2_X4 U_g25000 ( .A1(g24013), .A2(g24038), .ZN(g25000) );
OR2_X4 U_g25183 ( .A1(g24958), .A2(g24893), .ZN(g25183) );
OR2_X4 U_g25186 ( .A1(g24969), .A2(g24916), .ZN(g25186) );
OR2_X4 U_g25190 ( .A1(g24982), .A2(g24933), .ZN(g25190) );
OR2_X4 U_g25195 ( .A1(g24993), .A2(g24945), .ZN(g25195) );
OR2_X4 U_g25489 ( .A1(g24795), .A2(g16466), .ZN(g25489) );
OR2_X4 U_g25490 ( .A1(g24759), .A2(g23146), .ZN(g25490) );
OR2_X4 U_g25520 ( .A1(g24813), .A2(g23145), .ZN(g25520) );
OR2_X4 U_g25566 ( .A1(g24843), .A2(g23143), .ZN(g25566) );
OR2_X4 U_g26320 ( .A1(g25852), .A2(g25870), .ZN(g26320) );
OR2_X4 U_g26367 ( .A1(g25873), .A2(g25882), .ZN(g26367) );
OR2_X4 U_g26410 ( .A1(g25885), .A2(g25887), .ZN(g26410) );
OR2_X4 U_g26451 ( .A1(g25890), .A2(g25892), .ZN(g26451) );
OR2_X4 U_g26974 ( .A1(g26157), .A2(g23147), .ZN(g26974) );
OR3_X4 U_g27113 ( .A1(g1248), .A2(g1245), .A3(g26534), .ZN(g27113) );
OR2_X4 U_g28501 ( .A1(g27738), .A2(g25764), .ZN(g28501) );
OR2_X4 U_g28512 ( .A1(g26481), .A2(g27738), .ZN(g28512) );
OR2_X4 U_g28529 ( .A1(g27743), .A2(g25818), .ZN(g28529) );
OR2_X4 U_g28540 ( .A1(g26497), .A2(g27743), .ZN(g28540) );
OR2_X4 U_g28556 ( .A1(g27751), .A2(g25853), .ZN(g28556) );
OR2_X4 U_g28567 ( .A1(g26512), .A2(g27751), .ZN(g28567) );
OR2_X4 U_g28584 ( .A1(g27756), .A2(g25874), .ZN(g28584) );
OR2_X4 U_g28595 ( .A1(g26520), .A2(g27756), .ZN(g28595) );
OR3_X4 U_g29348 ( .A1(g1942), .A2(g1939), .A3(g29113), .ZN(g29348) );
OR3_X4 U_g30305 ( .A1(g2636), .A2(g2633), .A3(g30072), .ZN(g30305) );
NAND2_X4 U_I15167 ( .A1(g2981), .A2(g2874), .ZN(I15167) );
NAND2_X4 U_I15168 ( .A1(g2981), .A2(I15167), .ZN(I15168) );
NAND2_X4 U_I15169 ( .A1(g2874), .A2(I15167), .ZN(I15169) );
NAND2_X4 U_g7855 ( .A1(I15168), .A2(I15169), .ZN(g7855) );
NAND2_X4 U_I15183 ( .A1(g2975), .A2(g2978), .ZN(I15183) );
NAND2_X4 U_I15184 ( .A1(g2975), .A2(I15183), .ZN(I15184) );
NAND2_X4 U_I15185 ( .A1(g2978), .A2(I15183), .ZN(I15185) );
NAND2_X4 U_g7875 ( .A1(I15184), .A2(I15185), .ZN(g7875) );
NAND2_X4 U_I15190 ( .A1(g2956), .A2(g2959), .ZN(I15190) );
NAND2_X4 U_I15191 ( .A1(g2956), .A2(I15190), .ZN(I15191) );
NAND2_X4 U_I15192 ( .A1(g2959), .A2(I15190), .ZN(I15192) );
NAND2_X4 U_g7876 ( .A1(I15191), .A2(I15192), .ZN(g7876) );
NAND2_X4 U_I15204 ( .A1(g2969), .A2(g2972), .ZN(I15204) );
NAND2_X4 U_I15205 ( .A1(g2969), .A2(I15204), .ZN(I15205) );
NAND2_X4 U_I15206 ( .A1(g2972), .A2(I15204), .ZN(I15206) );
NAND2_X4 U_g7895 ( .A1(I15205), .A2(I15206), .ZN(g7895) );
NAND2_X4 U_I15211 ( .A1(g2947), .A2(g2953), .ZN(I15211) );
NAND2_X4 U_I15212 ( .A1(g2947), .A2(I15211), .ZN(I15212) );
NAND2_X4 U_I15213 ( .A1(g2953), .A2(I15211), .ZN(I15213) );
NAND2_X4 U_g7896 ( .A1(I15212), .A2(I15213), .ZN(g7896) );
NAND2_X4 U_I15237 ( .A1(g2963), .A2(g2966), .ZN(I15237) );
NAND2_X4 U_I15238 ( .A1(g2963), .A2(I15237), .ZN(I15238) );
NAND2_X4 U_I15239 ( .A1(g2966), .A2(I15237), .ZN(I15239) );
NAND2_X4 U_g7922 ( .A1(I15238), .A2(I15239), .ZN(g7922) );
NAND2_X4 U_I15244 ( .A1(g2941), .A2(g2944), .ZN(I15244) );
NAND2_X4 U_I15245 ( .A1(g2941), .A2(I15244), .ZN(I15245) );
NAND2_X4 U_I15246 ( .A1(g2944), .A2(I15244), .ZN(I15246) );
NAND2_X4 U_g7923 ( .A1(I15245), .A2(I15246), .ZN(g7923) );
NAND2_X4 U_I15276 ( .A1(g2935), .A2(g2938), .ZN(I15276) );
NAND2_X4 U_I15277 ( .A1(g2935), .A2(I15276), .ZN(I15277) );
NAND2_X4 U_I15278 ( .A1(g2938), .A2(I15276), .ZN(I15278) );
NAND2_X4 U_g7970 ( .A1(I15277), .A2(I15278), .ZN(g7970) );
NAND4_X4 U_g8381 ( .A1(g8182), .A2(g8120), .A3(g8044), .A4(g7989), .ZN(g8381) );
NAND2_X4 U_g8533 ( .A1(g3398), .A2(g3366), .ZN(g8533) );
NAND2_X4 U_g8547 ( .A1(g3398), .A2(g3366), .ZN(g8547) );
NAND2_X4 U_g8550 ( .A1(g3554), .A2(g3522), .ZN(g8550) );
NAND2_X4 U_g8560 ( .A1(g3554), .A2(g3522), .ZN(g8560) );
NAND2_X4 U_g8563 ( .A1(g3710), .A2(g3678), .ZN(g8563) );
NAND2_X4 U_g8571 ( .A1(g3710), .A2(g3678), .ZN(g8571) );
NAND2_X4 U_g8574 ( .A1(g3866), .A2(g3834), .ZN(g8574) );
NAND2_X4 U_g8577 ( .A1(g3866), .A2(g3834), .ZN(g8577) );
NAND2_X4 U_I16879 ( .A1(g4203), .A2(g3998), .ZN(I16879) );
NAND2_X4 U_I16880 ( .A1(g4203), .A2(I16879), .ZN(I16880) );
NAND2_X4 U_I16881 ( .A1(g3998), .A2(I16879), .ZN(I16881) );
NAND2_X4 U_g9883 ( .A1(I16880), .A2(I16881), .ZN(g9883) );
NAND2_X4 U_I16965 ( .A1(g4734), .A2(g4452), .ZN(I16965) );
NAND2_X4 U_I16966 ( .A1(g4734), .A2(I16965), .ZN(I16966) );
NAND2_X4 U_I16967 ( .A1(g4452), .A2(I16965), .ZN(I16967) );
NAND2_X4 U_g10003 ( .A1(I16966), .A2(I16967), .ZN(g10003) );
NAND2_X4 U_g10038 ( .A1(g7772), .A2(g3366), .ZN(g10038) );
NAND2_X4 U_I17059 ( .A1(g6637), .A2(g6309), .ZN(I17059) );
NAND2_X4 U_I17060 ( .A1(g6637), .A2(I17059), .ZN(I17060) );
NAND2_X4 U_I17061 ( .A1(g6309), .A2(I17059), .ZN(I17061) );
NAND2_X4 U_g10095 ( .A1(I17060), .A2(I17061), .ZN(g10095) );
NAND2_X4 U_g10147 ( .A1(g7788), .A2(g3522), .ZN(g10147) );
NAND2_X4 U_I17149 ( .A1(g7465), .A2(g7142), .ZN(I17149) );
NAND2_X4 U_I17150 ( .A1(g7465), .A2(I17149), .ZN(I17150) );
NAND2_X4 U_I17151 ( .A1(g7142), .A2(I17149), .ZN(I17151) );
NAND2_X4 U_g10185 ( .A1(I17150), .A2(I17151), .ZN(g10185) );
NAND2_X4 U_g10252 ( .A1(g7802), .A2(g3678), .ZN(g10252) );
NAND2_X4 U_g10354 ( .A1(g7815), .A2(g3834), .ZN(g10354) );
NAND2_X4 U_g10649 ( .A1(g3398), .A2(g6912), .ZN(g10649) );
NAND2_X4 U_g10676 ( .A1(g3398), .A2(g6678), .ZN(g10676) );
NAND2_X4 U_g10677 ( .A1(g3398), .A2(g6912), .ZN(g10677) );
NAND2_X4 U_g10679 ( .A1(g3554), .A2(g7162), .ZN(g10679) );
NAND2_X4 U_g10703 ( .A1(g3398), .A2(g6678), .ZN(g10703) );
NAND2_X4 U_g10705 ( .A1(g3554), .A2(g6980), .ZN(g10705) );
NAND2_X4 U_g10706 ( .A1(g3554), .A2(g7162), .ZN(g10706) );
NAND2_X4 U_g10708 ( .A1(g3710), .A2(g7358), .ZN(g10708) );
NAND2_X4 U_g10723 ( .A1(g3554), .A2(g6980), .ZN(g10723) );
NAND2_X4 U_g10725 ( .A1(g3710), .A2(g7230), .ZN(g10725) );
NAND2_X4 U_g10726 ( .A1(g3710), .A2(g7358), .ZN(g10726) );
NAND2_X4 U_g10728 ( .A1(g3866), .A2(g7488), .ZN(g10728) );
NAND2_X4 U_g10744 ( .A1(g3710), .A2(g7230), .ZN(g10744) );
NAND2_X4 U_g10746 ( .A1(g3866), .A2(g7426), .ZN(g10746) );
NAND2_X4 U_g10747 ( .A1(g3866), .A2(g7488), .ZN(g10747) );
NAND2_X4 U_g10763 ( .A1(g3866), .A2(g7426), .ZN(g10763) );
NAND2_X4 U_I18106 ( .A1(g7875), .A2(g7855), .ZN(I18106) );
NAND2_X4 U_I18107 ( .A1(g7875), .A2(I18106), .ZN(I18107) );
NAND2_X4 U_I18108 ( .A1(g7855), .A2(I18106), .ZN(I18108) );
NAND2_X4 U_g11188 ( .A1(I18107), .A2(I18108), .ZN(g11188) );
NAND2_X4 U_I18113 ( .A1(g3997), .A2(g8181), .ZN(I18113) );
NAND2_X4 U_I18114 ( .A1(g3997), .A2(I18113), .ZN(I18114) );
NAND2_X4 U_I18115 ( .A1(g8181), .A2(I18113), .ZN(I18115) );
NAND2_X4 U_g11189 ( .A1(I18114), .A2(I18115), .ZN(g11189) );
NAND2_X4 U_I18190 ( .A1(g7922), .A2(g7895), .ZN(I18190) );
NAND2_X4 U_I18191 ( .A1(g7922), .A2(I18190), .ZN(I18191) );
NAND2_X4 U_I18192 ( .A1(g7895), .A2(I18190), .ZN(I18192) );
NAND2_X4 U_g11262 ( .A1(I18191), .A2(I18192), .ZN(g11262) );
NAND2_X4 U_I18197 ( .A1(g7896), .A2(g7876), .ZN(I18197) );
NAND2_X4 U_I18198 ( .A1(g7896), .A2(I18197), .ZN(I18198) );
NAND2_X4 U_I18199 ( .A1(g7876), .A2(I18197), .ZN(I18199) );
NAND2_X4 U_g11263 ( .A1(I18198), .A2(I18199), .ZN(g11263) );
NAND2_X4 U_I18204 ( .A1(g7975), .A2(g4202), .ZN(I18204) );
NAND2_X4 U_I18205 ( .A1(g7975), .A2(I18204), .ZN(I18205) );
NAND2_X4 U_I18206 ( .A1(g4202), .A2(I18204), .ZN(I18206) );
NAND2_X4 U_g11264 ( .A1(I18205), .A2(I18206), .ZN(g11264) );
NAND2_X4 U_I18280 ( .A1(g7970), .A2(g7923), .ZN(I18280) );
NAND2_X4 U_I18281 ( .A1(g7970), .A2(I18280), .ZN(I18281) );
NAND2_X4 U_I18282 ( .A1(g7923), .A2(I18280), .ZN(I18282) );
NAND2_X4 U_g11330 ( .A1(I18281), .A2(I18282), .ZN(g11330) );
NAND2_X4 U_I18287 ( .A1(g8256), .A2(g8102), .ZN(I18287) );
NAND2_X4 U_I18288 ( .A1(g8256), .A2(I18287), .ZN(I18288) );
NAND2_X4 U_I18289 ( .A1(g8102), .A2(I18287), .ZN(I18289) );
NAND2_X4 U_g11331 ( .A1(I18288), .A2(I18289), .ZN(g11331) );
NAND2_X4 U_I18368 ( .A1(g4325), .A2(g4093), .ZN(I18368) );
NAND2_X4 U_I18369 ( .A1(g4325), .A2(I18368), .ZN(I18369) );
NAND2_X4 U_I18370 ( .A1(g4093), .A2(I18368), .ZN(I18370) );
NAND2_X4 U_g11410 ( .A1(I18369), .A2(I18370), .ZN(g11410) );
NAND2_X4 U_g11617 ( .A1(g8313), .A2(g2883), .ZN(g11617) );
NAND2_X4 U_I18799 ( .A1(g11410), .A2(g11331), .ZN(I18799) );
NAND2_X4 U_I18800 ( .A1(g11410), .A2(I18799), .ZN(I18800) );
NAND2_X4 U_I18801 ( .A1(g11331), .A2(I18799), .ZN(I18801) );
NAND2_X4 U_g11621 ( .A1(I18800), .A2(I18801), .ZN(g11621) );
NAND2_X4 U_g11661 ( .A1(g9534), .A2(g3366), .ZN(g11661) );
NAND2_X4 U_g11662 ( .A1(g9534), .A2(g3366), .ZN(g11662) );
NAND2_X4 U_g11672 ( .A1(g9534), .A2(g3366), .ZN(g11672) );
NAND2_X4 U_g11673 ( .A1(g9676), .A2(g3522), .ZN(g11673) );
NAND2_X4 U_g11674 ( .A1(g9676), .A2(g3522), .ZN(g11674) );
NAND2_X4 U_g11683 ( .A1(g9534), .A2(g3366), .ZN(g11683) );
NAND2_X4 U_g11684 ( .A1(g9676), .A2(g3522), .ZN(g11684) );
NAND2_X4 U_g11685 ( .A1(g9822), .A2(g3678), .ZN(g11685) );
NAND2_X4 U_g11686 ( .A1(g9822), .A2(g3678), .ZN(g11686) );
NAND2_X4 U_g11691 ( .A1(g9534), .A2(g3366), .ZN(g11691) );
NAND2_X4 U_g11692 ( .A1(g9676), .A2(g3522), .ZN(g11692) );
NAND2_X4 U_g11693 ( .A1(g9822), .A2(g3678), .ZN(g11693) );
NAND2_X4 U_g11694 ( .A1(g9968), .A2(g3834), .ZN(g11694) );
NAND2_X4 U_g11695 ( .A1(g9968), .A2(g3834), .ZN(g11695) );
NAND2_X4 U_g11696 ( .A1(g9534), .A2(g3366), .ZN(g11696) );
NAND2_X4 U_g11698 ( .A1(g9676), .A2(g3522), .ZN(g11698) );
NAND2_X4 U_g11699 ( .A1(g9822), .A2(g3678), .ZN(g11699) );
NAND2_X4 U_g11700 ( .A1(g9968), .A2(g3834), .ZN(g11700) );
NAND2_X4 U_g11701 ( .A1(g9534), .A2(g3366), .ZN(g11701) );
NAND2_X4 U_g11702 ( .A1(g9676), .A2(g3522), .ZN(g11702) );
NAND2_X4 U_g11704 ( .A1(g9822), .A2(g3678), .ZN(g11704) );
NAND2_X4 U_g11705 ( .A1(g9968), .A2(g3834), .ZN(g11705) );
NAND2_X4 U_g11707 ( .A1(g9534), .A2(g3366), .ZN(g11707) );
NAND2_X4 U_g11708 ( .A1(g9534), .A2(g3366), .ZN(g11708) );
NAND2_X4 U_g11709 ( .A1(g9676), .A2(g3522), .ZN(g11709) );
NAND2_X4 U_g11710 ( .A1(g9822), .A2(g3678), .ZN(g11710) );
NAND2_X4 U_g11712 ( .A1(g9968), .A2(g3834), .ZN(g11712) );
NAND2_X4 U_g11713 ( .A1(g10481), .A2(g9144), .ZN(g11713) );
NAND2_X4 U_g11716 ( .A1(g9534), .A2(g3366), .ZN(g11716) );
NAND2_X4 U_g11717 ( .A1(g9676), .A2(g3522), .ZN(g11717) );
NAND2_X4 U_g11718 ( .A1(g9676), .A2(g3522), .ZN(g11718) );
NAND2_X4 U_g11719 ( .A1(g9822), .A2(g3678), .ZN(g11719) );
NAND2_X4 U_g11720 ( .A1(g9968), .A2(g3834), .ZN(g11720) );
NAND2_X4 U_g11721 ( .A1(g9534), .A2(g3366), .ZN(g11721) );
NAND2_X4 U_g11722 ( .A1(g9676), .A2(g3522), .ZN(g11722) );
NAND2_X4 U_g11723 ( .A1(g9822), .A2(g3678), .ZN(g11723) );
NAND2_X4 U_g11724 ( .A1(g9822), .A2(g3678), .ZN(g11724) );
NAND2_X4 U_g11725 ( .A1(g9968), .A2(g3834), .ZN(g11725) );
NAND2_X4 U_g11726 ( .A1(g9676), .A2(g3522), .ZN(g11726) );
NAND2_X4 U_g11727 ( .A1(g9822), .A2(g3678), .ZN(g11727) );
NAND2_X4 U_g11728 ( .A1(g9968), .A2(g3834), .ZN(g11728) );
NAND2_X4 U_g11729 ( .A1(g9968), .A2(g3834), .ZN(g11729) );
NAND2_X4 U_g11730 ( .A1(g9822), .A2(g3678), .ZN(g11730) );
NAND2_X4 U_g11731 ( .A1(g9968), .A2(g3834), .ZN(g11731) );
NAND2_X4 U_g11733 ( .A1(g9968), .A2(g3834), .ZN(g11733) );
NAND2_X4 U_g12433 ( .A1(g2879), .A2(g10778), .ZN(g12433) );
NAND2_X4 U_g12486 ( .A1(g8278), .A2(g6448), .ZN(g12486) );
NAND2_X4 U_g12503 ( .A1(g8278), .A2(g5438), .ZN(g12503) );
NAND2_X4 U_g12506 ( .A1(g8287), .A2(g6713), .ZN(g12506) );
NAND2_X4 U_g12520 ( .A1(g8287), .A2(g5473), .ZN(g12520) );
NAND2_X4 U_g12523 ( .A1(g8296), .A2(g7015), .ZN(g12523) );
NAND2_X4 U_g12535 ( .A1(g8296), .A2(g5512), .ZN(g12535) );
NAND2_X4 U_g12538 ( .A1(g8305), .A2(g7265), .ZN(g12538) );
NAND2_X4 U_g12544 ( .A1(g8305), .A2(g5556), .ZN(g12544) );
NAND2_X4 U_I20031 ( .A1(g10003), .A2(g9883), .ZN(I20031) );
NAND2_X4 U_I20032 ( .A1(g10003), .A2(I20031), .ZN(I20032) );
NAND2_X4 U_I20033 ( .A1(g9883), .A2(I20031), .ZN(I20033) );
NAND2_X4 U_g12988 ( .A1(I20032), .A2(I20033), .ZN(g12988) );
NAND2_X4 U_I20048 ( .A1(g10185), .A2(g10095), .ZN(I20048) );
NAND2_X4 U_I20049 ( .A1(g10185), .A2(I20048), .ZN(I20049) );
NAND2_X4 U_I20050 ( .A1(g10095), .A2(I20048), .ZN(I20050) );
NAND2_X4 U_g12999 ( .A1(I20049), .A2(I20050), .ZN(g12999) );
NAND2_X4 U_g13020 ( .A1(g9534), .A2(g6912), .ZN(g13020) );
NAND2_X4 U_g13021 ( .A1(g9534), .A2(g6912), .ZN(g13021) );
NAND2_X4 U_g13026 ( .A1(g9534), .A2(g6678), .ZN(g13026) );
NAND2_X4 U_g13027 ( .A1(g9534), .A2(g6912), .ZN(g13027) );
NAND2_X4 U_g13028 ( .A1(g9534), .A2(g6678), .ZN(g13028) );
NAND2_X4 U_g13029 ( .A1(g9676), .A2(g7162), .ZN(g13029) );
NAND2_X4 U_g13030 ( .A1(g9676), .A2(g7162), .ZN(g13030) );
NAND2_X4 U_g13034 ( .A1(g9534), .A2(g6678), .ZN(g13034) );
NAND2_X4 U_g13035 ( .A1(g9534), .A2(g6912), .ZN(g13035) );
NAND2_X4 U_g13037 ( .A1(g9676), .A2(g6980), .ZN(g13037) );
NAND2_X4 U_g13038 ( .A1(g9676), .A2(g7162), .ZN(g13038) );
NAND2_X4 U_g13039 ( .A1(g9676), .A2(g6980), .ZN(g13039) );
NAND2_X4 U_g13040 ( .A1(g9822), .A2(g7358), .ZN(g13040) );
NAND2_X4 U_g13041 ( .A1(g9822), .A2(g7358), .ZN(g13041) );
NAND2_X4 U_g13044 ( .A1(g9534), .A2(g6678), .ZN(g13044) );
NAND2_X4 U_g13045 ( .A1(g9534), .A2(g6912), .ZN(g13045) );
NAND2_X4 U_g13047 ( .A1(g9676), .A2(g6980), .ZN(g13047) );
NAND2_X4 U_g13048 ( .A1(g9676), .A2(g7162), .ZN(g13048) );
NAND2_X4 U_g13050 ( .A1(g9822), .A2(g7230), .ZN(g13050) );
NAND2_X4 U_g13051 ( .A1(g9822), .A2(g7358), .ZN(g13051) );
NAND2_X4 U_g13052 ( .A1(g9822), .A2(g7230), .ZN(g13052) );
NAND2_X4 U_g13053 ( .A1(g9968), .A2(g7488), .ZN(g13053) );
NAND2_X4 U_g13054 ( .A1(g9968), .A2(g7488), .ZN(g13054) );
NAND2_X4 U_g13058 ( .A1(g9534), .A2(g6678), .ZN(g13058) );
NAND2_X4 U_g13059 ( .A1(g9534), .A2(g6912), .ZN(g13059) );
NAND2_X4 U_g13061 ( .A1(g9676), .A2(g6980), .ZN(g13061) );
NAND2_X4 U_g13062 ( .A1(g9676), .A2(g7162), .ZN(g13062) );
NAND2_X4 U_g13064 ( .A1(g9822), .A2(g7230), .ZN(g13064) );
NAND2_X4 U_g13065 ( .A1(g9822), .A2(g7358), .ZN(g13065) );
NAND2_X4 U_g13067 ( .A1(g9968), .A2(g7426), .ZN(g13067) );
NAND2_X4 U_g13068 ( .A1(g9968), .A2(g7488), .ZN(g13068) );
NAND2_X4 U_g13069 ( .A1(g9968), .A2(g7426), .ZN(g13069) );
NAND2_X4 U_g13071 ( .A1(g9534), .A2(g6678), .ZN(g13071) );
NAND2_X4 U_g13072 ( .A1(g9534), .A2(g6912), .ZN(g13072) );
NAND2_X4 U_g13074 ( .A1(g9676), .A2(g6980), .ZN(g13074) );
NAND2_X4 U_g13075 ( .A1(g9676), .A2(g7162), .ZN(g13075) );
NAND2_X4 U_g13077 ( .A1(g9822), .A2(g7230), .ZN(g13077) );
NAND2_X4 U_g13078 ( .A1(g9822), .A2(g7358), .ZN(g13078) );
NAND2_X4 U_g13080 ( .A1(g9968), .A2(g7426), .ZN(g13080) );
NAND2_X4 U_g13081 ( .A1(g9968), .A2(g7488), .ZN(g13081) );
NAND2_X4 U_g13087 ( .A1(g9534), .A2(g6678), .ZN(g13087) );
NAND2_X4 U_g13088 ( .A1(g9534), .A2(g6912), .ZN(g13088) );
NAND2_X4 U_g13089 ( .A1(g9534), .A2(g6912), .ZN(g13089) );
NAND2_X4 U_g13090 ( .A1(g9676), .A2(g6980), .ZN(g13090) );
NAND2_X4 U_g13091 ( .A1(g9676), .A2(g7162), .ZN(g13091) );
NAND2_X4 U_g13093 ( .A1(g9822), .A2(g7230), .ZN(g13093) );
NAND2_X4 U_g13094 ( .A1(g9822), .A2(g7358), .ZN(g13094) );
NAND2_X4 U_g13096 ( .A1(g9968), .A2(g7426), .ZN(g13096) );
NAND2_X4 U_g13097 ( .A1(g9968), .A2(g7488), .ZN(g13097) );
NAND2_X4 U_g13098 ( .A1(g9534), .A2(g6678), .ZN(g13098) );
NAND2_X4 U_g13099 ( .A1(g9534), .A2(g6912), .ZN(g13099) );
NAND2_X4 U_g13100 ( .A1(g9534), .A2(g6678), .ZN(g13100) );
NAND2_X4 U_g13102 ( .A1(g9676), .A2(g6980), .ZN(g13102) );
NAND2_X4 U_g13103 ( .A1(g9676), .A2(g7162), .ZN(g13103) );
NAND2_X4 U_g13104 ( .A1(g9676), .A2(g7162), .ZN(g13104) );
NAND2_X4 U_g13105 ( .A1(g9822), .A2(g7230), .ZN(g13105) );
NAND2_X4 U_g13106 ( .A1(g9822), .A2(g7358), .ZN(g13106) );
NAND2_X4 U_g13108 ( .A1(g9968), .A2(g7426), .ZN(g13108) );
NAND2_X4 U_g13109 ( .A1(g9968), .A2(g7488), .ZN(g13109) );
NAND2_X4 U_g13112 ( .A1(g9534), .A2(g6678), .ZN(g13112) );
NAND2_X4 U_g13113 ( .A1(g9534), .A2(g6912), .ZN(g13113) );
NAND2_X4 U_g13114 ( .A1(g9676), .A2(g6980), .ZN(g13114) );
NAND2_X4 U_g13115 ( .A1(g9676), .A2(g7162), .ZN(g13115) );
NAND2_X4 U_g13116 ( .A1(g9676), .A2(g6980), .ZN(g13116) );
NAND2_X4 U_g13118 ( .A1(g9822), .A2(g7230), .ZN(g13118) );
NAND2_X4 U_g13119 ( .A1(g9822), .A2(g7358), .ZN(g13119) );
NAND2_X4 U_g13120 ( .A1(g9822), .A2(g7358), .ZN(g13120) );
NAND2_X4 U_g13121 ( .A1(g9968), .A2(g7426), .ZN(g13121) );
NAND2_X4 U_g13122 ( .A1(g9968), .A2(g7488), .ZN(g13122) );
NAND2_X4 U_g13123 ( .A1(g9534), .A2(g6678), .ZN(g13123) );
NAND2_X4 U_g13125 ( .A1(g9676), .A2(g6980), .ZN(g13125) );
NAND2_X4 U_g13126 ( .A1(g9676), .A2(g7162), .ZN(g13126) );
NAND2_X4 U_g13127 ( .A1(g9822), .A2(g7230), .ZN(g13127) );
NAND2_X4 U_g13128 ( .A1(g9822), .A2(g7358), .ZN(g13128) );
NAND2_X4 U_g13129 ( .A1(g9822), .A2(g7230), .ZN(g13129) );
NAND2_X4 U_g13131 ( .A1(g9968), .A2(g7426), .ZN(g13131) );
NAND2_X4 U_g13132 ( .A1(g9968), .A2(g7488), .ZN(g13132) );
NAND2_X4 U_g13133 ( .A1(g9968), .A2(g7488), .ZN(g13133) );
NAND2_X4 U_g13134 ( .A1(g9676), .A2(g6980), .ZN(g13134) );
NAND2_X4 U_g13136 ( .A1(g9822), .A2(g7230), .ZN(g13136) );
NAND2_X4 U_g13137 ( .A1(g9822), .A2(g7358), .ZN(g13137) );
NAND2_X4 U_g13138 ( .A1(g9968), .A2(g7426), .ZN(g13138) );
NAND2_X4 U_g13139 ( .A1(g9968), .A2(g7488), .ZN(g13139) );
NAND2_X4 U_g13140 ( .A1(g9968), .A2(g7426), .ZN(g13140) );
NAND2_X4 U_g13142 ( .A1(g9822), .A2(g7230), .ZN(g13142) );
NAND2_X4 U_g13144 ( .A1(g9968), .A2(g7426), .ZN(g13144) );
NAND2_X4 U_g13145 ( .A1(g9968), .A2(g7488), .ZN(g13145) );
NAND2_X4 U_g13146 ( .A1(g9968), .A2(g7426), .ZN(g13146) );
NAND2_X4 U_g13147 ( .A1(g8278), .A2(g3306), .ZN(g13147) );
NAND2_X4 U_g13150 ( .A1(g8287), .A2(g3462), .ZN(g13150) );
NAND2_X4 U_g13156 ( .A1(g8296), .A2(g3618), .ZN(g13156) );
NAND2_X4 U_g13165 ( .A1(g8305), .A2(g3774), .ZN(g13165) );
NAND2_X4 U_g13245 ( .A1(g10779), .A2(g7901), .ZN(g13245) );
NAND2_X4 U_g13305 ( .A1(g8317), .A2(g2993), .ZN(g13305) );
NAND2_X4 U_I20429 ( .A1(g11262), .A2(g11188), .ZN(I20429) );
NAND2_X4 U_I20430 ( .A1(g11262), .A2(I20429), .ZN(I20430) );
NAND2_X4 U_I20431 ( .A1(g11188), .A2(I20429), .ZN(I20431) );
NAND2_X4 U_g13348 ( .A1(I20430), .A2(I20431), .ZN(g13348) );
NAND2_X4 U_I20465 ( .A1(g11330), .A2(g11263), .ZN(I20465) );
NAND2_X4 U_I20466 ( .A1(g11330), .A2(I20465), .ZN(I20466) );
NAND2_X4 U_I20467 ( .A1(g11263), .A2(I20465), .ZN(I20467) );
NAND2_X4 U_g13370 ( .A1(I20466), .A2(I20467), .ZN(g13370) );
NAND2_X4 U_I20504 ( .A1(g11264), .A2(g11189), .ZN(I20504) );
NAND2_X4 U_I20505 ( .A1(g11264), .A2(I20504), .ZN(I20505) );
NAND2_X4 U_I20506 ( .A1(g11189), .A2(I20504), .ZN(I20506) );
NAND2_X4 U_g13399 ( .A1(I20505), .A2(I20506), .ZN(g13399) );
NAND2_X4 U_g13476 ( .A1(g12565), .A2(g3254), .ZN(g13476) );
NAND2_X4 U_g13478 ( .A1(g12611), .A2(g3410), .ZN(g13478) );
NAND2_X4 U_g13482 ( .A1(g12657), .A2(g3566), .ZN(g13482) );
NAND2_X4 U_g13494 ( .A1(g12565), .A2(g3254), .ZN(g13494) );
NAND2_X4 U_g13495 ( .A1(g12611), .A2(g3410), .ZN(g13495) );
NAND2_X4 U_g13497 ( .A1(g12657), .A2(g3566), .ZN(g13497) );
NAND2_X4 U_g13501 ( .A1(g12711), .A2(g3722), .ZN(g13501) );
NAND2_X4 U_I20743 ( .A1(g11621), .A2(g13399), .ZN(I20743) );
NAND2_X4 U_I20744 ( .A1(g11621), .A2(I20743), .ZN(I20744) );
NAND2_X4 U_I20745 ( .A1(g13399), .A2(I20743), .ZN(I20745) );
NAND2_X4 U_g13507 ( .A1(I20744), .A2(I20745), .ZN(g13507) );
NAND2_X4 U_g13510 ( .A1(g12565), .A2(g3254), .ZN(g13510) );
NAND2_X4 U_g13511 ( .A1(g12611), .A2(g3410), .ZN(g13511) );
NAND2_X4 U_g13512 ( .A1(g12657), .A2(g3566), .ZN(g13512) );
NAND2_X4 U_g13514 ( .A1(g12711), .A2(g3722), .ZN(g13514) );
NAND2_X4 U_g13518 ( .A1(g12565), .A2(g3254), .ZN(g13518) );
NAND2_X4 U_g13524 ( .A1(g12611), .A2(g3410), .ZN(g13524) );
NAND2_X4 U_g13525 ( .A1(g12657), .A2(g3566), .ZN(g13525) );
NAND2_X4 U_g13526 ( .A1(g12711), .A2(g3722), .ZN(g13526) );
NAND2_X4 U_g13528 ( .A1(g12565), .A2(g3254), .ZN(g13528) );
NAND2_X4 U_g13529 ( .A1(g12611), .A2(g3410), .ZN(g13529) );
NAND2_X4 U_g13535 ( .A1(g12657), .A2(g3566), .ZN(g13535) );
NAND2_X4 U_g13536 ( .A1(g12711), .A2(g3722), .ZN(g13536) );
NAND2_X4 U_g13537 ( .A1(g12565), .A2(g3254), .ZN(g13537) );
NAND2_X4 U_g13538 ( .A1(g12565), .A2(g3254), .ZN(g13538) );
NAND2_X4 U_g13539 ( .A1(g12611), .A2(g3410), .ZN(g13539) );
NAND2_X4 U_g13540 ( .A1(g12657), .A2(g3566), .ZN(g13540) );
NAND2_X4 U_g13546 ( .A1(g12711), .A2(g3722), .ZN(g13546) );
NAND2_X4 U_g13547 ( .A1(g12565), .A2(g3254), .ZN(g13547) );
NAND2_X4 U_g13548 ( .A1(g12611), .A2(g3410), .ZN(g13548) );
NAND2_X4 U_g13549 ( .A1(g12611), .A2(g3410), .ZN(g13549) );
NAND2_X4 U_g13550 ( .A1(g12657), .A2(g3566), .ZN(g13550) );
NAND2_X4 U_g13551 ( .A1(g12711), .A2(g3722), .ZN(g13551) );
NAND2_X4 U_g13557 ( .A1(g12611), .A2(g3410), .ZN(g13557) );
NAND2_X4 U_g13558 ( .A1(g12657), .A2(g3566), .ZN(g13558) );
NAND2_X4 U_g13559 ( .A1(g12657), .A2(g3566), .ZN(g13559) );
NAND2_X4 U_g13560 ( .A1(g12711), .A2(g3722), .ZN(g13560) );
NAND2_X4 U_g13561 ( .A1(g12657), .A2(g3566), .ZN(g13561) );
NAND2_X4 U_g13562 ( .A1(g12711), .A2(g3722), .ZN(g13562) );
NAND2_X4 U_g13563 ( .A1(g12711), .A2(g3722), .ZN(g13563) );
NAND2_X4 U_g13564 ( .A1(g12711), .A2(g3722), .ZN(g13564) );
NAND2_X4 U_g13599 ( .A1(g12886), .A2(g3366), .ZN(g13599) );
NAND2_X4 U_g13611 ( .A1(g12926), .A2(g3522), .ZN(g13611) );
NAND2_X4 U_g13621 ( .A1(g12955), .A2(g3678), .ZN(g13621) );
NAND2_X4 U_g13633 ( .A1(g12984), .A2(g3834), .ZN(g13633) );
NAND2_X4 U_g13893 ( .A1(g8580), .A2(g12463), .ZN(g13893) );
NAND3_X4 U_g13915 ( .A1(g8822), .A2(g12473), .A3(g12463), .ZN(g13915) );
NAND2_X4 U_g13934 ( .A1(g8587), .A2(g12478), .ZN(g13934) );
NAND2_X4 U_g13957 ( .A1(g10730), .A2(g12473), .ZN(g13957) );
NAND3_X4 U_g13971 ( .A1(g8846), .A2(g12490), .A3(g12478), .ZN(g13971) );
NAND2_X4 U_g13990 ( .A1(g8594), .A2(g12495), .ZN(g13990) );
NAND2_X4 U_g14027 ( .A1(g10749), .A2(g12490), .ZN(g14027) );
NAND3_X4 U_g14041 ( .A1(g8873), .A2(g12510), .A3(g12495), .ZN(g14041) );
NAND2_X4 U_g14060 ( .A1(g8605), .A2(g12515), .ZN(g14060) );
NAND2_X4 U_g14118 ( .A1(g10767), .A2(g12510), .ZN(g14118) );
NAND3_X4 U_g14132 ( .A1(g8911), .A2(g12527), .A3(g12515), .ZN(g14132) );
NAND2_X4 U_g14233 ( .A1(g10773), .A2(g12527), .ZN(g14233) );
NAND3_X4 U_g15454 ( .A1(g9232), .A2(g9150), .A3(g12780), .ZN(g15454) );
NAND3_X4 U_g15540 ( .A1(g9310), .A2(g9174), .A3(g12819), .ZN(g15540) );
NAND3_X4 U_g15618 ( .A1(g9391), .A2(g9216), .A3(g12857), .ZN(g15618) );
NAND2_X4 U_g15660 ( .A1(g13401), .A2(g12354), .ZN(g15660) );
NAND2_X4 U_g15664 ( .A1(g12565), .A2(g6314), .ZN(g15664) );
NAND3_X4 U_g15694 ( .A1(g9488), .A2(g9277), .A3(g12898), .ZN(g15694) );
NAND2_X4 U_g15718 ( .A1(g13286), .A2(g12354), .ZN(g15718) );
NAND2_X4 U_g15719 ( .A1(g13401), .A2(g12392), .ZN(g15719) );
NAND2_X4 U_g15720 ( .A1(g12565), .A2(g6232), .ZN(g15720) );
NAND2_X4 U_g15721 ( .A1(g12565), .A2(g6314), .ZN(g15721) );
NAND2_X4 U_g15723 ( .A1(g12611), .A2(g6519), .ZN(g15723) );
NAND2_X4 U_g15756 ( .A1(g13313), .A2(g12354), .ZN(g15756) );
NAND2_X4 U_g15757 ( .A1(g11622), .A2(g12392), .ZN(g15757) );
NAND2_X4 U_g15758 ( .A1(g12565), .A2(g6232), .ZN(g15758) );
NAND2_X4 U_g15759 ( .A1(g12565), .A2(g6314), .ZN(g15759) );
NAND2_X4 U_g15760 ( .A1(g12611), .A2(g6369), .ZN(g15760) );
NAND2_X4 U_g15761 ( .A1(g12611), .A2(g6519), .ZN(g15761) );
NAND2_X4 U_g15763 ( .A1(g12657), .A2(g6783), .ZN(g15763) );
NAND2_X4 U_g15782 ( .A1(g13332), .A2(g12354), .ZN(g15782) );
NAND2_X4 U_g15783 ( .A1(g11643), .A2(g12392), .ZN(g15783) );
NAND2_X4 U_g15784 ( .A1(g12565), .A2(g6232), .ZN(g15784) );
NAND2_X4 U_g15785 ( .A1(g12565), .A2(g6314), .ZN(g15785) );
NAND2_X4 U_g15786 ( .A1(g12611), .A2(g6369), .ZN(g15786) );
NAND2_X4 U_g15787 ( .A1(g12611), .A2(g6519), .ZN(g15787) );
NAND2_X4 U_g15788 ( .A1(g12657), .A2(g6574), .ZN(g15788) );
NAND2_X4 U_g15789 ( .A1(g12657), .A2(g6783), .ZN(g15789) );
NAND2_X4 U_g15791 ( .A1(g12711), .A2(g7085), .ZN(g15791) );
NAND2_X4 U_g15803 ( .A1(g13375), .A2(g12354), .ZN(g15803) );
NAND2_X4 U_g15804 ( .A1(g11660), .A2(g12392), .ZN(g15804) );
NAND2_X4 U_g15805 ( .A1(g12565), .A2(g6232), .ZN(g15805) );
NAND2_X4 U_g15806 ( .A1(g12565), .A2(g6314), .ZN(g15806) );
NAND2_X4 U_g15807 ( .A1(g12611), .A2(g6369), .ZN(g15807) );
NAND2_X4 U_g15808 ( .A1(g12611), .A2(g6519), .ZN(g15808) );
NAND2_X4 U_g15809 ( .A1(g12657), .A2(g6574), .ZN(g15809) );
NAND2_X4 U_g15810 ( .A1(g12657), .A2(g6783), .ZN(g15810) );
NAND2_X4 U_g15811 ( .A1(g12711), .A2(g6838), .ZN(g15811) );
NAND2_X4 U_g15812 ( .A1(g12711), .A2(g7085), .ZN(g15812) );
NAND2_X4 U_I22062 ( .A1(g12999), .A2(g12988), .ZN(I22062) );
NAND2_X4 U_I22063 ( .A1(g12999), .A2(I22062), .ZN(I22063) );
NAND2_X4 U_I22064 ( .A1(g12988), .A2(I22062), .ZN(I22064) );
NAND2_X4 U_g15814 ( .A1(I22063), .A2(I22064), .ZN(g15814) );
NAND2_X4 U_g15818 ( .A1(g13024), .A2(g12354), .ZN(g15818) );
NAND2_X4 U_g15819 ( .A1(g13286), .A2(g12392), .ZN(g15819) );
NAND2_X4 U_g15820 ( .A1(g12565), .A2(g6232), .ZN(g15820) );
NAND2_X4 U_g15821 ( .A1(g12565), .A2(g6314), .ZN(g15821) );
NAND2_X4 U_g15822 ( .A1(g12611), .A2(g6369), .ZN(g15822) );
NAND2_X4 U_g15823 ( .A1(g12611), .A2(g6519), .ZN(g15823) );
NAND2_X4 U_g15824 ( .A1(g12657), .A2(g6574), .ZN(g15824) );
NAND2_X4 U_g15825 ( .A1(g12657), .A2(g6783), .ZN(g15825) );
NAND2_X4 U_g15826 ( .A1(g12711), .A2(g6838), .ZN(g15826) );
NAND2_X4 U_g15827 ( .A1(g12711), .A2(g7085), .ZN(g15827) );
NAND2_X4 U_g15830 ( .A1(g13310), .A2(g12392), .ZN(g15830) );
NAND2_X4 U_g15831 ( .A1(g13313), .A2(g12392), .ZN(g15831) );
NAND2_X4 U_g15832 ( .A1(g12565), .A2(g6232), .ZN(g15832) );
NAND2_X4 U_g15833 ( .A1(g12565), .A2(g6314), .ZN(g15833) );
NAND2_X4 U_g15834 ( .A1(g12611), .A2(g6369), .ZN(g15834) );
NAND2_X4 U_g15835 ( .A1(g12611), .A2(g6519), .ZN(g15835) );
NAND2_X4 U_g15836 ( .A1(g12657), .A2(g6574), .ZN(g15836) );
NAND2_X4 U_g15837 ( .A1(g12657), .A2(g6783), .ZN(g15837) );
NAND2_X4 U_g15838 ( .A1(g12711), .A2(g6838), .ZN(g15838) );
NAND2_X4 U_g15839 ( .A1(g12711), .A2(g7085), .ZN(g15839) );
NAND2_X4 U_g15841 ( .A1(g13331), .A2(g12392), .ZN(g15841) );
NAND2_X4 U_g15842 ( .A1(g13332), .A2(g12392), .ZN(g15842) );
NAND2_X4 U_g15843 ( .A1(g12565), .A2(g6314), .ZN(g15843) );
NAND2_X4 U_g15844 ( .A1(g12565), .A2(g6232), .ZN(g15844) );
NAND2_X4 U_g15845 ( .A1(g12565), .A2(g6314), .ZN(g15845) );
NAND2_X4 U_g15846 ( .A1(g12611), .A2(g6369), .ZN(g15846) );
NAND2_X4 U_g15847 ( .A1(g12611), .A2(g6519), .ZN(g15847) );
NAND2_X4 U_g15848 ( .A1(g12657), .A2(g6574), .ZN(g15848) );
NAND2_X4 U_g15849 ( .A1(g12657), .A2(g6783), .ZN(g15849) );
NAND2_X4 U_g15850 ( .A1(g12711), .A2(g6838), .ZN(g15850) );
NAND2_X4 U_g15851 ( .A1(g12711), .A2(g7085), .ZN(g15851) );
NAND2_X4 U_g15853 ( .A1(g13310), .A2(g12354), .ZN(g15853) );
NAND2_X4 U_g15854 ( .A1(g13353), .A2(g12392), .ZN(g15854) );
NAND2_X4 U_g15855 ( .A1(g13354), .A2(g12392), .ZN(g15855) );
NAND2_X4 U_g15856 ( .A1(g12565), .A2(g6232), .ZN(g15856) );
NAND2_X4 U_g15857 ( .A1(g12565), .A2(g6314), .ZN(g15857) );
NAND2_X4 U_g15858 ( .A1(g12565), .A2(g6232), .ZN(g15858) );
NAND2_X4 U_g15866 ( .A1(g12611), .A2(g6519), .ZN(g15866) );
NAND2_X4 U_g15867 ( .A1(g12611), .A2(g6369), .ZN(g15867) );
NAND2_X4 U_g15868 ( .A1(g12611), .A2(g6519), .ZN(g15868) );
NAND2_X4 U_g15869 ( .A1(g12657), .A2(g6574), .ZN(g15869) );
NAND2_X4 U_g15870 ( .A1(g12657), .A2(g6783), .ZN(g15870) );
NAND2_X4 U_g15871 ( .A1(g12711), .A2(g6838), .ZN(g15871) );
NAND2_X4 U_g15872 ( .A1(g12711), .A2(g7085), .ZN(g15872) );
NAND2_X4 U_g15877 ( .A1(g13374), .A2(g12392), .ZN(g15877) );
NAND2_X4 U_g15878 ( .A1(g13375), .A2(g12392), .ZN(g15878) );
NAND2_X4 U_g15879 ( .A1(g12565), .A2(g6232), .ZN(g15879) );
NAND2_X4 U_g15887 ( .A1(g12611), .A2(g6369), .ZN(g15887) );
NAND2_X4 U_g15888 ( .A1(g12611), .A2(g6519), .ZN(g15888) );
NAND2_X4 U_g15889 ( .A1(g12611), .A2(g6369), .ZN(g15889) );
NAND2_X4 U_g15897 ( .A1(g12657), .A2(g6783), .ZN(g15897) );
NAND2_X4 U_g15898 ( .A1(g12657), .A2(g6574), .ZN(g15898) );
NAND2_X4 U_g15899 ( .A1(g12657), .A2(g6783), .ZN(g15899) );
NAND2_X4 U_g15900 ( .A1(g12711), .A2(g6838), .ZN(g15900) );
NAND2_X4 U_g15901 ( .A1(g12711), .A2(g7085), .ZN(g15901) );
NAND2_X4 U_g15903 ( .A1(g13404), .A2(g12392), .ZN(g15903) );
NAND2_X4 U_g15912 ( .A1(g12611), .A2(g6369), .ZN(g15912) );
NAND2_X4 U_g15920 ( .A1(g12657), .A2(g6574), .ZN(g15920) );
NAND2_X4 U_g15921 ( .A1(g12657), .A2(g6783), .ZN(g15921) );
NAND2_X4 U_g15922 ( .A1(g12657), .A2(g6574), .ZN(g15922) );
NAND2_X4 U_g15930 ( .A1(g12711), .A2(g7085), .ZN(g15930) );
NAND2_X4 U_g15931 ( .A1(g12711), .A2(g6838), .ZN(g15931) );
NAND2_X4 U_g15932 ( .A1(g12711), .A2(g7085), .ZN(g15932) );
NAND2_X4 U_g15941 ( .A1(g12657), .A2(g6574), .ZN(g15941) );
NAND2_X4 U_g15949 ( .A1(g12711), .A2(g6838), .ZN(g15949) );
NAND2_X4 U_g15950 ( .A1(g12711), .A2(g7085), .ZN(g15950) );
NAND2_X4 U_g15951 ( .A1(g12711), .A2(g6838), .ZN(g15951) );
NAND2_X4 U_g15970 ( .A1(g12711), .A2(g6838), .ZN(g15970) );
NAND2_X4 U_g15990 ( .A1(g12886), .A2(g6912), .ZN(g15990) );
NAND2_X4 U_g15992 ( .A1(g12886), .A2(g6678), .ZN(g15992) );
NAND2_X4 U_g15993 ( .A1(g12926), .A2(g7162), .ZN(g15993) );
NAND2_X4 U_g15995 ( .A1(g12926), .A2(g6980), .ZN(g15995) );
NAND2_X4 U_g15996 ( .A1(g12955), .A2(g7358), .ZN(g15996) );
NAND2_X4 U_g15999 ( .A1(g12955), .A2(g7230), .ZN(g15999) );
NAND2_X4 U_g16000 ( .A1(g12984), .A2(g7488), .ZN(g16000) );
NAND2_X4 U_g16006 ( .A1(g12984), .A2(g7426), .ZN(g16006) );
NAND2_X4 U_g16085 ( .A1(g12883), .A2(g633), .ZN(g16085) );
NAND2_X4 U_g16123 ( .A1(g12923), .A2(g1319), .ZN(g16123) );
NAND2_X4 U_I22282 ( .A1(g2962), .A2(g13348), .ZN(I22282) );
NAND2_X4 U_I22283 ( .A1(g2962), .A2(I22282), .ZN(I22283) );
NAND2_X4 U_I22284 ( .A1(g13348), .A2(I22282), .ZN(I22284) );
NAND2_X4 U_g16132 ( .A1(I22283), .A2(I22284), .ZN(g16132) );
NAND2_X4 U_g16174 ( .A1(g12952), .A2(g2013), .ZN(g16174) );
NAND2_X4 U_I22316 ( .A1(g2934), .A2(g13370), .ZN(I22316) );
NAND2_X4 U_I22317 ( .A1(g2934), .A2(I22316), .ZN(I22317) );
NAND2_X4 U_I22318 ( .A1(g13370), .A2(I22316), .ZN(I22318) );
NAND2_X4 U_g16181 ( .A1(I22317), .A2(I22318), .ZN(g16181) );
NAND2_X4 U_g16233 ( .A1(g12981), .A2(g2707), .ZN(g16233) );
NAND2_X4 U_g16341 ( .A1(g12377), .A2(g12407), .ZN(g16341) );
NAND2_X4 U_g16412 ( .A1(g12565), .A2(g3254), .ZN(g16412) );
NAND2_X4 U_g16439 ( .A1(g13082), .A2(g2912), .ZN(g16439) );
NAND2_X4 U_g16442 ( .A1(g12565), .A2(g3254), .ZN(g16442) );
NAND2_X4 U_g16446 ( .A1(g12611), .A2(g3410), .ZN(g16446) );
NAND2_X4 U_g16463 ( .A1(g13004), .A2(g3018), .ZN(g16463) );
NAND2_X4 U_g16536 ( .A1(g15873), .A2(g2896), .ZN(g16536) );
NAND2_X4 U_I22630 ( .A1(g13507), .A2(g15978), .ZN(I22630) );
NAND2_X4 U_I22631 ( .A1(g13507), .A2(I22630), .ZN(I22631) );
NAND2_X4 U_I22632 ( .A1(g15978), .A2(I22630), .ZN(I22632) );
NAND2_X4 U_g16566 ( .A1(I22631), .A2(I22632), .ZN(g16566) );
NAND2_X4 U_I22705 ( .A1(g13348), .A2(g15661), .ZN(I22705) );
NAND2_X4 U_I22706 ( .A1(g13348), .A2(I22705), .ZN(I22706) );
NAND2_X4 U_I22707 ( .A1(g15661), .A2(I22705), .ZN(I22707) );
NAND2_X4 U_g16662 ( .A1(I22706), .A2(I22707), .ZN(g16662) );
NAND2_X4 U_I22884 ( .A1(g13370), .A2(g15661), .ZN(I22884) );
NAND2_X4 U_I22885 ( .A1(g13370), .A2(I22884), .ZN(I22885) );
NAND2_X4 U_I22886 ( .A1(g15661), .A2(I22884), .ZN(I22886) );
NAND2_X4 U_g16935 ( .A1(I22885), .A2(I22886), .ZN(g16935) );
NAND2_X4 U_I22900 ( .A1(g15022), .A2(g14000), .ZN(I22900) );
NAND2_X4 U_I22901 ( .A1(g15022), .A2(I22900), .ZN(I22901) );
NAND2_X4 U_I22902 ( .A1(g14000), .A2(I22900), .ZN(I22902) );
NAND2_X4 U_g16965 ( .A1(I22901), .A2(I22902), .ZN(g16965) );
NAND2_X4 U_I22917 ( .A1(g15096), .A2(g13945), .ZN(I22917) );
NAND2_X4 U_I22918 ( .A1(g15096), .A2(I22917), .ZN(I22918) );
NAND2_X4 U_I22919 ( .A1(g13945), .A2(I22917), .ZN(I22919) );
NAND2_X4 U_g16985 ( .A1(I22918), .A2(I22919), .ZN(g16985) );
NAND2_X4 U_I22924 ( .A1(g15118), .A2(g14091), .ZN(I22924) );
NAND2_X4 U_I22925 ( .A1(g15118), .A2(I22924), .ZN(I22925) );
NAND2_X4 U_I22926 ( .A1(g14091), .A2(I22924), .ZN(I22926) );
NAND2_X4 U_g16986 ( .A1(I22925), .A2(I22926), .ZN(g16986) );
NAND2_X4 U_I22936 ( .A1(g9150), .A2(g13906), .ZN(I22936) );
NAND2_X4 U_I22937 ( .A1(g9150), .A2(I22936), .ZN(I22937) );
NAND2_X4 U_I22938 ( .A1(g13906), .A2(I22936), .ZN(I22938) );
NAND2_X4 U_g16992 ( .A1(I22937), .A2(I22938), .ZN(g16992) );
NAND2_X4 U_I22945 ( .A1(g15188), .A2(g14015), .ZN(I22945) );
NAND2_X4 U_I22946 ( .A1(g15188), .A2(I22945), .ZN(I22946) );
NAND2_X4 U_I22947 ( .A1(g14015), .A2(I22945), .ZN(I22947) );
NAND2_X4 U_g16995 ( .A1(I22946), .A2(I22947), .ZN(g16995) );
NAND2_X4 U_I22952 ( .A1(g15210), .A2(g14206), .ZN(I22952) );
NAND2_X4 U_I22953 ( .A1(g15210), .A2(I22952), .ZN(I22953) );
NAND2_X4 U_I22954 ( .A1(g14206), .A2(I22952), .ZN(I22954) );
NAND2_X4 U_g16996 ( .A1(I22953), .A2(I22954), .ZN(g16996) );
NAND2_X4 U_I22962 ( .A1(g9161), .A2(g13885), .ZN(I22962) );
NAND2_X4 U_I22963 ( .A1(g9161), .A2(I22962), .ZN(I22963) );
NAND2_X4 U_I22964 ( .A1(g13885), .A2(I22962), .ZN(I22964) );
NAND2_X4 U_g17000 ( .A1(I22963), .A2(I22964), .ZN(g17000) );
NAND2_X4 U_I22972 ( .A1(g9174), .A2(g13962), .ZN(I22972) );
NAND2_X4 U_I22973 ( .A1(g9174), .A2(I22972), .ZN(I22973) );
NAND2_X4 U_I22974 ( .A1(g13962), .A2(I22972), .ZN(I22974) );
NAND2_X4 U_g17016 ( .A1(I22973), .A2(I22974), .ZN(g17016) );
NAND2_X4 U_I22981 ( .A1(g15274), .A2(g14106), .ZN(I22981) );
NAND2_X4 U_I22982 ( .A1(g15274), .A2(I22981), .ZN(I22982) );
NAND2_X4 U_I22983 ( .A1(g14106), .A2(I22981), .ZN(I22983) );
NAND2_X4 U_g17019 ( .A1(I22982), .A2(I22983), .ZN(g17019) );
NAND2_X4 U_I22988 ( .A1(g15296), .A2(g14321), .ZN(I22988) );
NAND2_X4 U_I22989 ( .A1(g15296), .A2(I22988), .ZN(I22989) );
NAND2_X4 U_I22990 ( .A1(g14321), .A2(I22988), .ZN(I22990) );
NAND2_X4 U_g17020 ( .A1(I22989), .A2(I22990), .ZN(g17020) );
NAND2_X4 U_I22998 ( .A1(g9187), .A2(g13872), .ZN(I22998) );
NAND2_X4 U_I22999 ( .A1(g9187), .A2(I22998), .ZN(I22999) );
NAND2_X4 U_I23000 ( .A1(g13872), .A2(I22998), .ZN(I23000) );
NAND2_X4 U_g17024 ( .A1(I22999), .A2(I23000), .ZN(g17024) );
NAND2_X4 U_I23008 ( .A1(g9203), .A2(g13926), .ZN(I23008) );
NAND2_X4 U_I23009 ( .A1(g9203), .A2(I23008), .ZN(I23009) );
NAND2_X4 U_I23010 ( .A1(g13926), .A2(I23008), .ZN(I23010) );
NAND2_X4 U_g17030 ( .A1(I23009), .A2(I23010), .ZN(g17030) );
NAND2_X4 U_I23018 ( .A1(g9216), .A2(g14032), .ZN(I23018) );
NAND2_X4 U_I23019 ( .A1(g9216), .A2(I23018), .ZN(I23019) );
NAND2_X4 U_I23020 ( .A1(g14032), .A2(I23018), .ZN(I23020) );
NAND2_X4 U_g17046 ( .A1(I23019), .A2(I23020), .ZN(g17046) );
NAND2_X4 U_I23027 ( .A1(g15366), .A2(g14221), .ZN(I23027) );
NAND2_X4 U_I23028 ( .A1(g15366), .A2(I23027), .ZN(I23028) );
NAND2_X4 U_I23029 ( .A1(g14221), .A2(I23027), .ZN(I23029) );
NAND2_X4 U_g17049 ( .A1(I23028), .A2(I23029), .ZN(g17049) );
NAND2_X4 U_I23034 ( .A1(g9232), .A2(g13864), .ZN(I23034) );
NAND2_X4 U_I23035 ( .A1(g9232), .A2(I23034), .ZN(I23035) );
NAND2_X4 U_I23036 ( .A1(g13864), .A2(I23034), .ZN(I23036) );
NAND2_X4 U_g17050 ( .A1(I23035), .A2(I23036), .ZN(g17050) );
NAND2_X4 U_I23045 ( .A1(g9248), .A2(g13894), .ZN(I23045) );
NAND2_X4 U_I23046 ( .A1(g9248), .A2(I23045), .ZN(I23046) );
NAND2_X4 U_I23047 ( .A1(g13894), .A2(I23045), .ZN(I23047) );
NAND2_X4 U_g17058 ( .A1(I23046), .A2(I23047), .ZN(g17058) );
NAND2_X4 U_I23055 ( .A1(g9264), .A2(g13982), .ZN(I23055) );
NAND2_X4 U_I23056 ( .A1(g9264), .A2(I23055), .ZN(I23056) );
NAND2_X4 U_I23057 ( .A1(g13982), .A2(I23055), .ZN(I23057) );
NAND2_X4 U_g17064 ( .A1(I23056), .A2(I23057), .ZN(g17064) );
NAND2_X4 U_I23065 ( .A1(g9277), .A2(g14123), .ZN(I23065) );
NAND2_X4 U_I23066 ( .A1(g9277), .A2(I23065), .ZN(I23066) );
NAND2_X4 U_I23067 ( .A1(g14123), .A2(I23065), .ZN(I23067) );
NAND2_X4 U_g17080 ( .A1(I23066), .A2(I23067), .ZN(g17080) );
NAND2_X4 U_I23074 ( .A1(g9293), .A2(g13856), .ZN(I23074) );
NAND2_X4 U_I23075 ( .A1(g9293), .A2(I23074), .ZN(I23075) );
NAND2_X4 U_I23076 ( .A1(g13856), .A2(I23074), .ZN(I23076) );
NAND2_X4 U_g17083 ( .A1(I23075), .A2(I23076), .ZN(g17083) );
NAND2_X4 U_I23082 ( .A1(g9310), .A2(g13879), .ZN(I23082) );
NAND2_X4 U_I23083 ( .A1(g9310), .A2(I23082), .ZN(I23083) );
NAND2_X4 U_I23084 ( .A1(g13879), .A2(I23082), .ZN(I23084) );
NAND2_X4 U_g17085 ( .A1(I23083), .A2(I23084), .ZN(g17085) );
NAND2_X4 U_I23093 ( .A1(g9326), .A2(g13935), .ZN(I23093) );
NAND2_X4 U_I23094 ( .A1(g9326), .A2(I23093), .ZN(I23094) );
NAND2_X4 U_I23095 ( .A1(g13935), .A2(I23093), .ZN(I23095) );
NAND2_X4 U_g17093 ( .A1(I23094), .A2(I23095), .ZN(g17093) );
NAND2_X4 U_I23103 ( .A1(g9342), .A2(g14052), .ZN(I23103) );
NAND2_X4 U_I23104 ( .A1(g9342), .A2(I23103), .ZN(I23104) );
NAND2_X4 U_I23105 ( .A1(g14052), .A2(I23103), .ZN(I23105) );
NAND2_X4 U_g17099 ( .A1(I23104), .A2(I23105), .ZN(g17099) );
NAND2_X4 U_I23113 ( .A1(g9356), .A2(g13848), .ZN(I23113) );
NAND2_X4 U_I23114 ( .A1(g9356), .A2(I23113), .ZN(I23114) );
NAND2_X4 U_I23115 ( .A1(g13848), .A2(I23113), .ZN(I23115) );
NAND2_X4 U_g17115 ( .A1(I23114), .A2(I23115), .ZN(g17115) );
NAND2_X4 U_g17118 ( .A1(g13915), .A2(g13893), .ZN(g17118) );
NAND2_X4 U_I23123 ( .A1(g9374), .A2(g13866), .ZN(I23123) );
NAND2_X4 U_I23124 ( .A1(g9374), .A2(I23123), .ZN(I23124) );
NAND2_X4 U_I23125 ( .A1(g13866), .A2(I23123), .ZN(I23125) );
NAND2_X4 U_g17121 ( .A1(I23124), .A2(I23125), .ZN(g17121) );
NAND2_X4 U_I23131 ( .A1(g9391), .A2(g13901), .ZN(I23131) );
NAND2_X4 U_I23132 ( .A1(g9391), .A2(I23131), .ZN(I23132) );
NAND2_X4 U_I23133 ( .A1(g13901), .A2(I23131), .ZN(I23133) );
NAND2_X4 U_g17123 ( .A1(I23132), .A2(I23133), .ZN(g17123) );
NAND2_X4 U_I23142 ( .A1(g9407), .A2(g13991), .ZN(I23142) );
NAND2_X4 U_I23143 ( .A1(g9407), .A2(I23142), .ZN(I23143) );
NAND2_X4 U_I23144 ( .A1(g13991), .A2(I23142), .ZN(I23144) );
NAND2_X4 U_g17131 ( .A1(I23143), .A2(I23144), .ZN(g17131) );
NAND2_X4 U_I23152 ( .A1(g9427), .A2(g14061), .ZN(I23152) );
NAND2_X4 U_I23153 ( .A1(g9427), .A2(I23152), .ZN(I23153) );
NAND2_X4 U_I23154 ( .A1(g14061), .A2(I23152), .ZN(I23154) );
NAND2_X4 U_g17137 ( .A1(I23153), .A2(I23154), .ZN(g17137) );
NAND2_X4 U_g17139 ( .A1(g13957), .A2(g13915), .ZN(g17139) );
NAND2_X4 U_I23161 ( .A1(g9453), .A2(g13857), .ZN(I23161) );
NAND2_X4 U_I23162 ( .A1(g9453), .A2(I23161), .ZN(I23162) );
NAND2_X4 U_I23163 ( .A1(g13857), .A2(I23161), .ZN(I23163) );
NAND2_X4 U_g17142 ( .A1(I23162), .A2(I23163), .ZN(g17142) );
NAND2_X4 U_g17145 ( .A1(g13971), .A2(g13934), .ZN(g17145) );
NAND2_X4 U_I23171 ( .A1(g9471), .A2(g13881), .ZN(I23171) );
NAND2_X4 U_I23172 ( .A1(g9471), .A2(I23171), .ZN(I23172) );
NAND2_X4 U_I23173 ( .A1(g13881), .A2(I23171), .ZN(I23173) );
NAND2_X4 U_g17148 ( .A1(I23172), .A2(I23173), .ZN(g17148) );
NAND2_X4 U_I23179 ( .A1(g9488), .A2(g13942), .ZN(I23179) );
NAND2_X4 U_I23180 ( .A1(g9488), .A2(I23179), .ZN(I23180) );
NAND2_X4 U_I23181 ( .A1(g13942), .A2(I23179), .ZN(I23181) );
NAND2_X4 U_g17150 ( .A1(I23180), .A2(I23181), .ZN(g17150) );
NAND2_X4 U_I23190 ( .A1(g9507), .A2(g13999), .ZN(I23190) );
NAND2_X4 U_I23191 ( .A1(g9507), .A2(I23190), .ZN(I23191) );
NAND2_X4 U_I23192 ( .A1(g13999), .A2(I23190), .ZN(I23192) );
NAND2_X4 U_g17158 ( .A1(I23191), .A2(I23192), .ZN(g17158) );
NAND2_X4 U_g17159 ( .A1(g14642), .A2(g14657), .ZN(g17159) );
NAND2_X4 U_I23198 ( .A1(g9569), .A2(g14176), .ZN(I23198) );
NAND2_X4 U_I23199 ( .A1(g9569), .A2(I23198), .ZN(I23199) );
NAND2_X4 U_I23200 ( .A1(g14176), .A2(I23198), .ZN(I23200) );
NAND2_X4 U_g17160 ( .A1(I23199), .A2(I23200), .ZN(g17160) );
NAND2_X4 U_g17162 ( .A1(g14027), .A2(g13971), .ZN(g17162) );
NAND2_X4 U_I23207 ( .A1(g9595), .A2(g13867), .ZN(I23207) );
NAND2_X4 U_I23208 ( .A1(g9595), .A2(I23207), .ZN(I23208) );
NAND2_X4 U_I23209 ( .A1(g13867), .A2(I23207), .ZN(I23209) );
NAND2_X4 U_g17165 ( .A1(I23208), .A2(I23209), .ZN(g17165) );
NAND2_X4 U_g17168 ( .A1(g14041), .A2(g13990), .ZN(g17168) );
NAND2_X4 U_I23217 ( .A1(g9613), .A2(g13903), .ZN(I23217) );
NAND2_X4 U_I23218 ( .A1(g9613), .A2(I23217), .ZN(I23218) );
NAND2_X4 U_I23219 ( .A1(g13903), .A2(I23217), .ZN(I23219) );
NAND2_X4 U_g17171 ( .A1(I23218), .A2(I23219), .ZN(g17171) );
NAND2_X4 U_I23225 ( .A1(g9649), .A2(g14090), .ZN(I23225) );
NAND2_X4 U_I23226 ( .A1(g9649), .A2(I23225), .ZN(I23226) );
NAND2_X4 U_I23227 ( .A1(g14090), .A2(I23225), .ZN(I23227) );
NAND2_X4 U_g17173 ( .A1(I23226), .A2(I23227), .ZN(g17173) );
NAND2_X4 U_g17174 ( .A1(g14669), .A2(g14691), .ZN(g17174) );
NAND2_X4 U_I23233 ( .A1(g9711), .A2(g14291), .ZN(I23233) );
NAND2_X4 U_I23234 ( .A1(g9711), .A2(I23233), .ZN(I23234) );
NAND2_X4 U_I23235 ( .A1(g14291), .A2(I23233), .ZN(I23235) );
NAND2_X4 U_g17175 ( .A1(I23234), .A2(I23235), .ZN(g17175) );
NAND2_X4 U_g17177 ( .A1(g14118), .A2(g14041), .ZN(g17177) );
NAND2_X4 U_I23242 ( .A1(g9737), .A2(g13882), .ZN(I23242) );
NAND2_X4 U_I23243 ( .A1(g9737), .A2(I23242), .ZN(I23243) );
NAND2_X4 U_I23244 ( .A1(g13882), .A2(I23242), .ZN(I23244) );
NAND2_X4 U_g17180 ( .A1(I23243), .A2(I23244), .ZN(g17180) );
NAND2_X4 U_g17183 ( .A1(g14132), .A2(g14060), .ZN(g17183) );
NAND2_X4 U_I23256 ( .A1(g9795), .A2(g14205), .ZN(I23256) );
NAND2_X4 U_I23257 ( .A1(g9795), .A2(I23256), .ZN(I23257) );
NAND2_X4 U_I23258 ( .A1(g14205), .A2(I23256), .ZN(I23258) );
NAND2_X4 U_g17190 ( .A1(I23257), .A2(I23258), .ZN(g17190) );
NAND2_X4 U_g17191 ( .A1(g14703), .A2(g14725), .ZN(g17191) );
NAND2_X4 U_I23264 ( .A1(g9857), .A2(g14413), .ZN(I23264) );
NAND2_X4 U_I23265 ( .A1(g9857), .A2(I23264), .ZN(I23265) );
NAND2_X4 U_I23266 ( .A1(g14413), .A2(I23264), .ZN(I23266) );
NAND2_X4 U_g17192 ( .A1(I23265), .A2(I23266), .ZN(g17192) );
NAND2_X4 U_g17194 ( .A1(g14233), .A2(g14132), .ZN(g17194) );
NAND2_X4 U_I23277 ( .A1(g9941), .A2(g14320), .ZN(I23277) );
NAND2_X4 U_I23278 ( .A1(g9941), .A2(I23277), .ZN(I23278) );
NAND2_X4 U_I23279 ( .A1(g14320), .A2(I23277), .ZN(I23279) );
NAND2_X4 U_g17201 ( .A1(I23278), .A2(I23279), .ZN(g17201) );
NAND2_X4 U_g17202 ( .A1(g14737), .A2(g14753), .ZN(g17202) );
NAND2_X4 U_I23806 ( .A1(g14062), .A2(g9150), .ZN(I23806) );
NAND2_X4 U_I23807 ( .A1(g14062), .A2(I23806), .ZN(I23807) );
NAND2_X4 U_I23808 ( .A1(g9150), .A2(I23806), .ZN(I23808) );
NAND2_X4 U_g17729 ( .A1(I23807), .A2(I23808), .ZN(g17729) );
NAND2_X4 U_I23878 ( .A1(g14001), .A2(g9187), .ZN(I23878) );
NAND2_X4 U_I23879 ( .A1(g14001), .A2(I23878), .ZN(I23879) );
NAND2_X4 U_I23880 ( .A1(g9187), .A2(I23878), .ZN(I23880) );
NAND2_X4 U_g17807 ( .A1(I23879), .A2(I23880), .ZN(g17807) );
NAND2_X4 U_I23893 ( .A1(g14177), .A2(g9174), .ZN(I23893) );
NAND2_X4 U_I23894 ( .A1(g14177), .A2(I23893), .ZN(I23894) );
NAND2_X4 U_I23895 ( .A1(g9174), .A2(I23893), .ZN(I23895) );
NAND2_X4 U_g17830 ( .A1(I23894), .A2(I23895), .ZN(g17830) );
NAND2_X4 U_I23941 ( .A1(g13946), .A2(g9293), .ZN(I23941) );
NAND2_X4 U_I23942 ( .A1(g13946), .A2(I23941), .ZN(I23942) );
NAND2_X4 U_I23943 ( .A1(g9293), .A2(I23941), .ZN(I23943) );
NAND2_X4 U_g17887 ( .A1(I23942), .A2(I23943), .ZN(g17887) );
NAND2_X4 U_I23958 ( .A1(g6513), .A2(g14171), .ZN(I23958) );
NAND2_X4 U_I23959 ( .A1(g6513), .A2(I23958), .ZN(I23959) );
NAND2_X4 U_I23960 ( .A1(g14171), .A2(I23958), .ZN(I23960) );
NAND2_X4 U_g17913 ( .A1(I23959), .A2(I23960), .ZN(g17913) );
NAND2_X4 U_I23966 ( .A1(g14092), .A2(g9248), .ZN(I23966) );
NAND2_X4 U_I23967 ( .A1(g14092), .A2(I23966), .ZN(I23967) );
NAND2_X4 U_I23968 ( .A1(g9248), .A2(I23966), .ZN(I23968) );
NAND2_X4 U_g17919 ( .A1(I23967), .A2(I23968), .ZN(g17919) );
NAND2_X4 U_I23981 ( .A1(g14292), .A2(g9216), .ZN(I23981) );
NAND2_X4 U_I23982 ( .A1(g14292), .A2(I23981), .ZN(I23982) );
NAND2_X4 U_I23983 ( .A1(g9216), .A2(I23981), .ZN(I23983) );
NAND2_X4 U_g17942 ( .A1(I23982), .A2(I23983), .ZN(g17942) );
NAND2_X4 U_I24005 ( .A1(g7548), .A2(g15814), .ZN(I24005) );
NAND2_X4 U_I24006 ( .A1(g7548), .A2(I24005), .ZN(I24006) );
NAND2_X4 U_I24007 ( .A1(g15814), .A2(I24005), .ZN(I24007) );
NAND2_X4 U_g17968 ( .A1(I24006), .A2(I24007), .ZN(g17968) );
NAND2_X4 U_I24015 ( .A1(g13907), .A2(g9427), .ZN(I24015) );
NAND2_X4 U_I24016 ( .A1(g13907), .A2(I24015), .ZN(I24016) );
NAND2_X4 U_I24017 ( .A1(g9427), .A2(I24015), .ZN(I24017) );
NAND2_X4 U_g17979 ( .A1(I24016), .A2(I24017), .ZN(g17979) );
NAND2_X4 U_g17985 ( .A1(g14641), .A2(g9636), .ZN(g17985) );
NAND2_X4 U_I24028 ( .A1(g6201), .A2(g14086), .ZN(I24028) );
NAND2_X4 U_I24029 ( .A1(g6201), .A2(I24028), .ZN(I24029) );
NAND2_X4 U_I24030 ( .A1(g14086), .A2(I24028), .ZN(I24030) );
NAND2_X4 U_g17992 ( .A1(I24029), .A2(I24030), .ZN(g17992) );
NAND2_X4 U_I24036 ( .A1(g14016), .A2(g9374), .ZN(I24036) );
NAND2_X4 U_I24037 ( .A1(g14016), .A2(I24036), .ZN(I24037) );
NAND2_X4 U_I24038 ( .A1(g9374), .A2(I24036), .ZN(I24038) );
NAND2_X4 U_g17998 ( .A1(I24037), .A2(I24038), .ZN(g17998) );
NAND2_X4 U_I24053 ( .A1(g6777), .A2(g14286), .ZN(I24053) );
NAND2_X4 U_I24054 ( .A1(g6777), .A2(I24053), .ZN(I24054) );
NAND2_X4 U_I24055 ( .A1(g14286), .A2(I24053), .ZN(I24055) );
NAND2_X4 U_g18024 ( .A1(I24054), .A2(I24055), .ZN(g18024) );
NAND2_X4 U_I24061 ( .A1(g14207), .A2(g9326), .ZN(I24061) );
NAND2_X4 U_I24062 ( .A1(g14207), .A2(I24061), .ZN(I24062) );
NAND2_X4 U_I24063 ( .A1(g9326), .A2(I24061), .ZN(I24063) );
NAND2_X4 U_g18030 ( .A1(I24062), .A2(I24063), .ZN(g18030) );
NAND2_X4 U_I24076 ( .A1(g14414), .A2(g9277), .ZN(I24076) );
NAND2_X4 U_I24077 ( .A1(g14414), .A2(I24076), .ZN(I24077) );
NAND2_X4 U_I24078 ( .A1(g9277), .A2(I24076), .ZN(I24078) );
NAND2_X4 U_g18053 ( .A1(I24077), .A2(I24078), .ZN(g18053) );
NAND2_X4 U_I24091 ( .A1(g13886), .A2(g15096), .ZN(I24091) );
NAND2_X4 U_I24092 ( .A1(g13886), .A2(I24091), .ZN(I24092) );
NAND2_X4 U_I24093 ( .A1(g15096), .A2(I24091), .ZN(I24093) );
NAND2_X4 U_g18079 ( .A1(I24092), .A2(I24093), .ZN(g18079) );
NAND2_X4 U_I24102 ( .A1(g6363), .A2(g14011), .ZN(I24102) );
NAND2_X4 U_I24103 ( .A1(g6363), .A2(I24102), .ZN(I24103) );
NAND2_X4 U_I24104 ( .A1(g14011), .A2(I24102), .ZN(I24104) );
NAND2_X4 U_g18090 ( .A1(I24103), .A2(I24104), .ZN(g18090) );
NAND2_X4 U_I24110 ( .A1(g13963), .A2(g9569), .ZN(I24110) );
NAND2_X4 U_I24111 ( .A1(g13963), .A2(I24110), .ZN(I24111) );
NAND2_X4 U_I24112 ( .A1(g9569), .A2(I24110), .ZN(I24112) );
NAND2_X4 U_g18096 ( .A1(I24111), .A2(I24112), .ZN(g18096) );
NAND2_X4 U_g18102 ( .A1(g14668), .A2(g9782), .ZN(g18102) );
NAND2_X4 U_I24123 ( .A1(g6290), .A2(g14201), .ZN(I24123) );
NAND2_X4 U_I24124 ( .A1(g6290), .A2(I24123), .ZN(I24124) );
NAND2_X4 U_I24125 ( .A1(g14201), .A2(I24123), .ZN(I24125) );
NAND2_X4 U_g18109 ( .A1(I24124), .A2(I24125), .ZN(g18109) );
NAND2_X4 U_I24131 ( .A1(g14107), .A2(g9471), .ZN(I24131) );
NAND2_X4 U_I24132 ( .A1(g14107), .A2(I24131), .ZN(I24132) );
NAND2_X4 U_I24133 ( .A1(g9471), .A2(I24131), .ZN(I24133) );
NAND2_X4 U_g18115 ( .A1(I24132), .A2(I24133), .ZN(g18115) );
NAND2_X4 U_I24148 ( .A1(g7079), .A2(g14408), .ZN(I24148) );
NAND2_X4 U_I24149 ( .A1(g7079), .A2(I24148), .ZN(I24149) );
NAND2_X4 U_I24150 ( .A1(g14408), .A2(I24148), .ZN(I24150) );
NAND2_X4 U_g18141 ( .A1(I24149), .A2(I24150), .ZN(g18141) );
NAND2_X4 U_I24156 ( .A1(g14322), .A2(g9407), .ZN(I24156) );
NAND2_X4 U_I24157 ( .A1(g14322), .A2(I24156), .ZN(I24157) );
NAND2_X4 U_I24158 ( .A1(g9407), .A2(I24156), .ZN(I24158) );
NAND2_X4 U_g18147 ( .A1(I24157), .A2(I24158), .ZN(g18147) );
NAND2_X4 U_I24178 ( .A1(g13873), .A2(g9161), .ZN(I24178) );
NAND2_X4 U_I24179 ( .A1(g13873), .A2(I24178), .ZN(I24179) );
NAND2_X4 U_I24180 ( .A1(g9161), .A2(I24178), .ZN(I24180) );
NAND2_X4 U_g18183 ( .A1(I24179), .A2(I24180), .ZN(g18183) );
NAND2_X4 U_I24186 ( .A1(g6177), .A2(g13958), .ZN(I24186) );
NAND2_X4 U_I24187 ( .A1(g6177), .A2(I24186), .ZN(I24187) );
NAND2_X4 U_I24188 ( .A1(g13958), .A2(I24186), .ZN(I24188) );
NAND2_X4 U_g18189 ( .A1(I24187), .A2(I24188), .ZN(g18189) );
NAND2_X4 U_I24194 ( .A1(g13927), .A2(g15188), .ZN(I24194) );
NAND2_X4 U_I24195 ( .A1(g13927), .A2(I24194), .ZN(I24195) );
NAND2_X4 U_I24196 ( .A1(g15188), .A2(I24194), .ZN(I24196) );
NAND2_X4 U_g18195 ( .A1(I24195), .A2(I24196), .ZN(g18195) );
NAND2_X4 U_I24205 ( .A1(g6568), .A2(g14102), .ZN(I24205) );
NAND2_X4 U_I24206 ( .A1(g6568), .A2(I24205), .ZN(I24206) );
NAND2_X4 U_I24207 ( .A1(g14102), .A2(I24205), .ZN(I24207) );
NAND2_X4 U_g18206 ( .A1(I24206), .A2(I24207), .ZN(g18206) );
NAND2_X4 U_I24213 ( .A1(g14033), .A2(g9711), .ZN(I24213) );
NAND2_X4 U_I24214 ( .A1(g14033), .A2(I24213), .ZN(I24214) );
NAND2_X4 U_I24215 ( .A1(g9711), .A2(I24213), .ZN(I24215) );
NAND2_X4 U_g18212 ( .A1(I24214), .A2(I24215), .ZN(g18212) );
NAND2_X4 U_g18218 ( .A1(g14702), .A2(g9928), .ZN(g18218) );
NAND2_X4 U_I24226 ( .A1(g6427), .A2(g14316), .ZN(I24226) );
NAND2_X4 U_I24227 ( .A1(g6427), .A2(I24226), .ZN(I24227) );
NAND2_X4 U_I24228 ( .A1(g14316), .A2(I24226), .ZN(I24228) );
NAND2_X4 U_g18225 ( .A1(I24227), .A2(I24228), .ZN(g18225) );
NAND2_X4 U_I24234 ( .A1(g14222), .A2(g9613), .ZN(I24234) );
NAND2_X4 U_I24235 ( .A1(g14222), .A2(I24234), .ZN(I24235) );
NAND2_X4 U_I24236 ( .A1(g9613), .A2(I24234), .ZN(I24236) );
NAND2_X4 U_g18231 ( .A1(I24235), .A2(I24236), .ZN(g18231) );
NAND2_X4 U_I24251 ( .A1(g7329), .A2(g14520), .ZN(I24251) );
NAND2_X4 U_I24252 ( .A1(g7329), .A2(I24251), .ZN(I24252) );
NAND2_X4 U_I24253 ( .A1(g14520), .A2(I24251), .ZN(I24253) );
NAND2_X4 U_g18257 ( .A1(I24252), .A2(I24253), .ZN(g18257) );
NAND2_X4 U_I24263 ( .A1(g14342), .A2(g9232), .ZN(I24263) );
NAND2_X4 U_I24264 ( .A1(g14342), .A2(I24263), .ZN(I24264) );
NAND2_X4 U_I24265 ( .A1(g9232), .A2(I24263), .ZN(I24265) );
NAND2_X4 U_g18270 ( .A1(I24264), .A2(I24265), .ZN(g18270) );
NAND2_X4 U_I24271 ( .A1(g6180), .A2(g13922), .ZN(I24271) );
NAND2_X4 U_I24272 ( .A1(g6180), .A2(I24271), .ZN(I24272) );
NAND2_X4 U_I24273 ( .A1(g13922), .A2(I24271), .ZN(I24273) );
NAND2_X4 U_g18276 ( .A1(I24272), .A2(I24273), .ZN(g18276) );
NAND2_X4 U_I24278 ( .A1(g6284), .A2(g13918), .ZN(I24278) );
NAND2_X4 U_I24279 ( .A1(g6284), .A2(I24278), .ZN(I24279) );
NAND2_X4 U_I24280 ( .A1(g13918), .A2(I24278), .ZN(I24280) );
NAND2_X4 U_g18277 ( .A1(I24279), .A2(I24280), .ZN(g18277) );
NAND2_X4 U_I24290 ( .A1(g13895), .A2(g9203), .ZN(I24290) );
NAND2_X4 U_I24291 ( .A1(g13895), .A2(I24290), .ZN(I24291) );
NAND2_X4 U_I24292 ( .A1(g9203), .A2(I24290), .ZN(I24292) );
NAND2_X4 U_g18290 ( .A1(I24291), .A2(I24292), .ZN(g18290) );
NAND2_X4 U_I24298 ( .A1(g6209), .A2(g14028), .ZN(I24298) );
NAND2_X4 U_I24299 ( .A1(g6209), .A2(I24298), .ZN(I24299) );
NAND2_X4 U_I24300 ( .A1(g14028), .A2(I24298), .ZN(I24300) );
NAND2_X4 U_g18296 ( .A1(I24299), .A2(I24300), .ZN(g18296) );
NAND2_X4 U_I24306 ( .A1(g13983), .A2(g15274), .ZN(I24306) );
NAND2_X4 U_I24307 ( .A1(g13983), .A2(I24306), .ZN(I24307) );
NAND2_X4 U_I24308 ( .A1(g15274), .A2(I24306), .ZN(I24308) );
NAND2_X4 U_g18302 ( .A1(I24307), .A2(I24308), .ZN(g18302) );
NAND2_X4 U_I24317 ( .A1(g6832), .A2(g14217), .ZN(I24317) );
NAND2_X4 U_I24318 ( .A1(g6832), .A2(I24317), .ZN(I24318) );
NAND2_X4 U_I24319 ( .A1(g14217), .A2(I24317), .ZN(I24319) );
NAND2_X4 U_g18313 ( .A1(I24318), .A2(I24319), .ZN(g18313) );
NAND2_X4 U_I24325 ( .A1(g14124), .A2(g9857), .ZN(I24325) );
NAND2_X4 U_I24326 ( .A1(g14124), .A2(I24325), .ZN(I24326) );
NAND2_X4 U_I24327 ( .A1(g9857), .A2(I24325), .ZN(I24327) );
NAND2_X4 U_g18319 ( .A1(I24326), .A2(I24327), .ZN(g18319) );
NAND2_X4 U_g18325 ( .A1(g14736), .A2(g10082), .ZN(g18325) );
NAND2_X4 U_I24338 ( .A1(g6632), .A2(g14438), .ZN(I24338) );
NAND2_X4 U_I24339 ( .A1(g6632), .A2(I24338), .ZN(I24339) );
NAND2_X4 U_I24340 ( .A1(g14438), .A2(I24338), .ZN(I24340) );
NAND2_X4 U_g18332 ( .A1(I24339), .A2(I24340), .ZN(g18332) );
NAND2_X4 U_I24351 ( .A1(g14238), .A2(g9356), .ZN(I24351) );
NAND2_X4 U_I24352 ( .A1(g14238), .A2(I24351), .ZN(I24352) );
NAND2_X4 U_I24353 ( .A1(g9356), .A2(I24351), .ZN(I24353) );
NAND2_X4 U_g18346 ( .A1(I24352), .A2(I24353), .ZN(g18346) );
NAND2_X4 U_I24361 ( .A1(g6157), .A2(g14525), .ZN(I24361) );
NAND2_X4 U_I24362 ( .A1(g6157), .A2(I24361), .ZN(I24362) );
NAND2_X4 U_I24363 ( .A1(g14525), .A2(I24361), .ZN(I24363) );
NAND2_X4 U_g18354 ( .A1(I24362), .A2(I24363), .ZN(g18354) );
NAND2_X4 U_I24372 ( .A1(g14454), .A2(g9310), .ZN(I24372) );
NAND2_X4 U_I24373 ( .A1(g14454), .A2(I24372), .ZN(I24373) );
NAND2_X4 U_I24374 ( .A1(g9310), .A2(I24372), .ZN(I24374) );
NAND2_X4 U_g18363 ( .A1(I24373), .A2(I24374), .ZN(g18363) );
NAND2_X4 U_I24380 ( .A1(g6212), .A2(g13978), .ZN(I24380) );
NAND2_X4 U_I24381 ( .A1(g6212), .A2(I24380), .ZN(I24381) );
NAND2_X4 U_I24382 ( .A1(g13978), .A2(I24380), .ZN(I24382) );
NAND2_X4 U_g18369 ( .A1(I24381), .A2(I24382), .ZN(g18369) );
NAND2_X4 U_I24387 ( .A1(g6421), .A2(g13974), .ZN(I24387) );
NAND2_X4 U_I24388 ( .A1(g6421), .A2(I24387), .ZN(I24388) );
NAND2_X4 U_I24389 ( .A1(g13974), .A2(I24387), .ZN(I24389) );
NAND2_X4 U_g18370 ( .A1(I24388), .A2(I24389), .ZN(g18370) );
NAND2_X4 U_I24399 ( .A1(g13936), .A2(g9264), .ZN(I24399) );
NAND2_X4 U_I24400 ( .A1(g13936), .A2(I24399), .ZN(I24400) );
NAND2_X4 U_I24401 ( .A1(g9264), .A2(I24399), .ZN(I24401) );
NAND2_X4 U_g18383 ( .A1(I24400), .A2(I24401), .ZN(g18383) );
NAND2_X4 U_I24407 ( .A1(g6298), .A2(g14119), .ZN(I24407) );
NAND2_X4 U_I24408 ( .A1(g6298), .A2(I24407), .ZN(I24408) );
NAND2_X4 U_I24409 ( .A1(g14119), .A2(I24407), .ZN(I24409) );
NAND2_X4 U_g18389 ( .A1(I24408), .A2(I24409), .ZN(g18389) );
NAND2_X4 U_I24415 ( .A1(g14053), .A2(g15366), .ZN(I24415) );
NAND2_X4 U_I24416 ( .A1(g14053), .A2(I24415), .ZN(I24416) );
NAND2_X4 U_I24417 ( .A1(g15366), .A2(I24415), .ZN(I24417) );
NAND2_X4 U_g18395 ( .A1(I24416), .A2(I24417), .ZN(g18395) );
NAND2_X4 U_I24426 ( .A1(g7134), .A2(g14332), .ZN(I24426) );
NAND2_X4 U_I24427 ( .A1(g7134), .A2(I24426), .ZN(I24427) );
NAND2_X4 U_I24428 ( .A1(g14332), .A2(I24426), .ZN(I24428) );
NAND2_X4 U_g18406 ( .A1(I24427), .A2(I24428), .ZN(g18406) );
NAND2_X4 U_I24436 ( .A1(g14153), .A2(g15022), .ZN(I24436) );
NAND2_X4 U_I24437 ( .A1(g14153), .A2(I24436), .ZN(I24437) );
NAND2_X4 U_I24438 ( .A1(g15022), .A2(I24436), .ZN(I24438) );
NAND2_X4 U_g18419 ( .A1(I24437), .A2(I24438), .ZN(g18419) );
NAND2_X4 U_I24443 ( .A1(g14148), .A2(g9507), .ZN(I24443) );
NAND2_X4 U_I24444 ( .A1(g14148), .A2(I24443), .ZN(I24444) );
NAND2_X4 U_I24445 ( .A1(g9507), .A2(I24443), .ZN(I24445) );
NAND2_X4 U_g18424 ( .A1(I24444), .A2(I24445), .ZN(g18424) );
NAND2_X4 U_I24452 ( .A1(g6142), .A2(g14450), .ZN(I24452) );
NAND2_X4 U_I24453 ( .A1(g6142), .A2(I24452), .ZN(I24453) );
NAND2_X4 U_I24454 ( .A1(g14450), .A2(I24452), .ZN(I24454) );
NAND2_X4 U_g18431 ( .A1(I24453), .A2(I24454), .ZN(g18431) );
NAND2_X4 U_I24464 ( .A1(g14360), .A2(g9453), .ZN(I24464) );
NAND2_X4 U_I24465 ( .A1(g14360), .A2(I24464), .ZN(I24465) );
NAND2_X4 U_I24466 ( .A1(g9453), .A2(I24464), .ZN(I24466) );
NAND2_X4 U_g18441 ( .A1(I24465), .A2(I24466), .ZN(g18441) );
NAND2_X4 U_I24474 ( .A1(g6184), .A2(g14580), .ZN(I24474) );
NAND2_X4 U_I24475 ( .A1(g6184), .A2(I24474), .ZN(I24475) );
NAND2_X4 U_I24476 ( .A1(g14580), .A2(I24474), .ZN(I24476) );
NAND2_X4 U_g18449 ( .A1(I24475), .A2(I24476), .ZN(g18449) );
NAND2_X4 U_I24485 ( .A1(g14541), .A2(g9391), .ZN(I24485) );
NAND2_X4 U_I24486 ( .A1(g14541), .A2(I24485), .ZN(I24486) );
NAND2_X4 U_I24487 ( .A1(g9391), .A2(I24485), .ZN(I24487) );
NAND2_X4 U_g18458 ( .A1(I24486), .A2(I24487), .ZN(g18458) );
NAND2_X4 U_I24493 ( .A1(g6301), .A2(g14048), .ZN(I24493) );
NAND2_X4 U_I24494 ( .A1(g6301), .A2(I24493), .ZN(I24494) );
NAND2_X4 U_I24495 ( .A1(g14048), .A2(I24493), .ZN(I24495) );
NAND2_X4 U_g18464 ( .A1(I24494), .A2(I24495), .ZN(g18464) );
NAND2_X4 U_I24500 ( .A1(g6626), .A2(g14044), .ZN(I24500) );
NAND2_X4 U_I24501 ( .A1(g6626), .A2(I24500), .ZN(I24501) );
NAND2_X4 U_I24502 ( .A1(g14044), .A2(I24500), .ZN(I24502) );
NAND2_X4 U_g18465 ( .A1(I24501), .A2(I24502), .ZN(g18465) );
NAND2_X4 U_I24512 ( .A1(g13992), .A2(g9342), .ZN(I24512) );
NAND2_X4 U_I24513 ( .A1(g13992), .A2(I24512), .ZN(I24513) );
NAND2_X4 U_I24514 ( .A1(g9342), .A2(I24512), .ZN(I24514) );
NAND2_X4 U_g18478 ( .A1(I24513), .A2(I24514), .ZN(g18478) );
NAND2_X4 U_I24520 ( .A1(g6435), .A2(g14234), .ZN(I24520) );
NAND2_X4 U_I24521 ( .A1(g6435), .A2(I24520), .ZN(I24521) );
NAND2_X4 U_I24522 ( .A1(g14234), .A2(I24520), .ZN(I24522) );
NAND2_X4 U_g18484 ( .A1(I24521), .A2(I24522), .ZN(g18484) );
NAND2_X4 U_I24530 ( .A1(g6707), .A2(g14355), .ZN(I24530) );
NAND2_X4 U_I24531 ( .A1(g6707), .A2(I24530), .ZN(I24531) );
NAND2_X4 U_I24532 ( .A1(g14355), .A2(I24530), .ZN(I24532) );
NAND2_X4 U_g18491 ( .A1(I24531), .A2(I24532), .ZN(g18491) );
NAND2_X4 U_I24537 ( .A1(g14268), .A2(g15118), .ZN(I24537) );
NAND2_X4 U_I24538 ( .A1(g14268), .A2(I24537), .ZN(I24538) );
NAND2_X4 U_I24539 ( .A1(g15118), .A2(I24537), .ZN(I24539) );
NAND2_X4 U_g18492 ( .A1(I24538), .A2(I24539), .ZN(g18492) );
NAND2_X4 U_I24544 ( .A1(g14263), .A2(g9649), .ZN(I24544) );
NAND2_X4 U_I24545 ( .A1(g14263), .A2(I24544), .ZN(I24545) );
NAND2_X4 U_I24546 ( .A1(g9649), .A2(I24544), .ZN(I24546) );
NAND2_X4 U_g18497 ( .A1(I24545), .A2(I24546), .ZN(g18497) );
NAND2_X4 U_I24553 ( .A1(g6163), .A2(g14537), .ZN(I24553) );
NAND2_X4 U_I24554 ( .A1(g6163), .A2(I24553), .ZN(I24554) );
NAND2_X4 U_I24555 ( .A1(g14537), .A2(I24553), .ZN(I24555) );
NAND2_X4 U_g18504 ( .A1(I24554), .A2(I24555), .ZN(g18504) );
NAND2_X4 U_I24565 ( .A1(g14472), .A2(g9595), .ZN(I24565) );
NAND2_X4 U_I24566 ( .A1(g14472), .A2(I24565), .ZN(I24566) );
NAND2_X4 U_I24567 ( .A1(g9595), .A2(I24565), .ZN(I24567) );
NAND2_X4 U_g18514 ( .A1(I24566), .A2(I24567), .ZN(g18514) );
NAND2_X4 U_I24575 ( .A1(g6216), .A2(g14614), .ZN(I24575) );
NAND2_X4 U_I24576 ( .A1(g6216), .A2(I24575), .ZN(I24576) );
NAND2_X4 U_I24577 ( .A1(g14614), .A2(I24575), .ZN(I24577) );
NAND2_X4 U_g18522 ( .A1(I24576), .A2(I24577), .ZN(g18522) );
NAND2_X4 U_I24586 ( .A1(g14596), .A2(g9488), .ZN(I24586) );
NAND2_X4 U_I24587 ( .A1(g14596), .A2(I24586), .ZN(I24587) );
NAND2_X4 U_I24588 ( .A1(g9488), .A2(I24586), .ZN(I24588) );
NAND2_X4 U_g18531 ( .A1(I24587), .A2(I24588), .ZN(g18531) );
NAND2_X4 U_I24594 ( .A1(g6438), .A2(g14139), .ZN(I24594) );
NAND2_X4 U_I24595 ( .A1(g6438), .A2(I24594), .ZN(I24595) );
NAND2_X4 U_I24596 ( .A1(g14139), .A2(I24594), .ZN(I24596) );
NAND2_X4 U_g18537 ( .A1(I24595), .A2(I24596), .ZN(g18537) );
NAND2_X4 U_I24601 ( .A1(g6890), .A2(g14135), .ZN(I24601) );
NAND2_X4 U_I24602 ( .A1(g6890), .A2(I24601), .ZN(I24602) );
NAND2_X4 U_I24603 ( .A1(g14135), .A2(I24601), .ZN(I24603) );
NAND2_X4 U_g18538 ( .A1(I24602), .A2(I24603), .ZN(g18538) );
NAND2_X4 U_I24611 ( .A1(g15814), .A2(g15978), .ZN(I24611) );
NAND2_X4 U_I24612 ( .A1(g15814), .A2(I24611), .ZN(I24612) );
NAND2_X4 U_I24613 ( .A1(g15978), .A2(I24611), .ZN(I24613) );
NAND2_X4 U_g18542 ( .A1(I24612), .A2(I24613), .ZN(g18542) );
NAND2_X4 U_I24624 ( .A1(g6136), .A2(g14252), .ZN(I24624) );
NAND2_X4 U_I24625 ( .A1(g6136), .A2(I24624), .ZN(I24625) );
NAND2_X4 U_I24626 ( .A1(g14252), .A2(I24624), .ZN(I24626) );
NAND2_X4 U_g18553 ( .A1(I24625), .A2(I24626), .ZN(g18553) );
NAND2_X4 U_I24632 ( .A1(g7009), .A2(g14467), .ZN(I24632) );
NAND2_X4 U_I24633 ( .A1(g7009), .A2(I24632), .ZN(I24633) );
NAND2_X4 U_I24634 ( .A1(g14467), .A2(I24632), .ZN(I24634) );
NAND2_X4 U_g18555 ( .A1(I24633), .A2(I24634), .ZN(g18555) );
NAND2_X4 U_I24639 ( .A1(g14390), .A2(g15210), .ZN(I24639) );
NAND2_X4 U_I24640 ( .A1(g14390), .A2(I24639), .ZN(I24640) );
NAND2_X4 U_I24641 ( .A1(g15210), .A2(I24639), .ZN(I24641) );
NAND2_X4 U_g18556 ( .A1(I24640), .A2(I24641), .ZN(g18556) );
NAND2_X4 U_I24646 ( .A1(g14385), .A2(g9795), .ZN(I24646) );
NAND2_X4 U_I24647 ( .A1(g14385), .A2(I24646), .ZN(I24647) );
NAND2_X4 U_I24648 ( .A1(g9795), .A2(I24646), .ZN(I24648) );
NAND2_X4 U_g18561 ( .A1(I24647), .A2(I24648), .ZN(g18561) );
NAND2_X4 U_I24655 ( .A1(g6190), .A2(g14592), .ZN(I24655) );
NAND2_X4 U_I24656 ( .A1(g6190), .A2(I24655), .ZN(I24656) );
NAND2_X4 U_I24657 ( .A1(g14592), .A2(I24655), .ZN(I24657) );
NAND2_X4 U_g18568 ( .A1(I24656), .A2(I24657), .ZN(g18568) );
NAND2_X4 U_I24667 ( .A1(g14559), .A2(g9737), .ZN(I24667) );
NAND2_X4 U_I24668 ( .A1(g14559), .A2(I24667), .ZN(I24668) );
NAND2_X4 U_I24669 ( .A1(g9737), .A2(I24667), .ZN(I24669) );
NAND2_X4 U_g18578 ( .A1(I24668), .A2(I24669), .ZN(g18578) );
NAND2_X4 U_I24677 ( .A1(g6305), .A2(g14637), .ZN(I24677) );
NAND2_X4 U_I24678 ( .A1(g6305), .A2(I24677), .ZN(I24678) );
NAND2_X4 U_I24679 ( .A1(g14637), .A2(I24677), .ZN(I24679) );
NAND2_X4 U_g18586 ( .A1(I24678), .A2(I24679), .ZN(g18586) );
NAND2_X4 U_I24694 ( .A1(g6146), .A2(g14374), .ZN(I24694) );
NAND2_X4 U_I24695 ( .A1(g6146), .A2(I24694), .ZN(I24695) );
NAND2_X4 U_I24696 ( .A1(g14374), .A2(I24694), .ZN(I24696) );
NAND2_X4 U_g18603 ( .A1(I24695), .A2(I24696), .ZN(g18603) );
NAND2_X4 U_I24702 ( .A1(g7259), .A2(g14554), .ZN(I24702) );
NAND2_X4 U_I24703 ( .A1(g7259), .A2(I24702), .ZN(I24703) );
NAND2_X4 U_I24704 ( .A1(g14554), .A2(I24702), .ZN(I24704) );
NAND2_X4 U_g18605 ( .A1(I24703), .A2(I24704), .ZN(g18605) );
NAND2_X4 U_I24709 ( .A1(g14502), .A2(g15296), .ZN(I24709) );
NAND2_X4 U_I24710 ( .A1(g14502), .A2(I24709), .ZN(I24710) );
NAND2_X4 U_I24711 ( .A1(g15296), .A2(I24709), .ZN(I24711) );
NAND2_X4 U_g18606 ( .A1(I24710), .A2(I24711), .ZN(g18606) );
NAND2_X4 U_I24716 ( .A1(g14497), .A2(g9941), .ZN(I24716) );
NAND2_X4 U_I24717 ( .A1(g14497), .A2(I24716), .ZN(I24717) );
NAND2_X4 U_I24718 ( .A1(g9941), .A2(I24716), .ZN(I24718) );
NAND2_X4 U_g18611 ( .A1(I24717), .A2(I24718), .ZN(g18611) );
NAND2_X4 U_I24725 ( .A1(g6222), .A2(g14626), .ZN(I24725) );
NAND2_X4 U_I24726 ( .A1(g6222), .A2(I24725), .ZN(I24726) );
NAND2_X4 U_I24727 ( .A1(g14626), .A2(I24725), .ZN(I24727) );
NAND2_X4 U_g18618 ( .A1(I24726), .A2(I24727), .ZN(g18618) );
NAND2_X4 U_I24743 ( .A1(g6167), .A2(g14486), .ZN(I24743) );
NAND2_X4 U_I24744 ( .A1(g6167), .A2(I24743), .ZN(I24744) );
NAND2_X4 U_I24745 ( .A1(g14486), .A2(I24743), .ZN(I24745) );
NAND2_X4 U_g18635 ( .A1(I24744), .A2(I24745), .ZN(g18635) );
NAND2_X4 U_I24751 ( .A1(g7455), .A2(g14609), .ZN(I24751) );
NAND2_X4 U_I24752 ( .A1(g7455), .A2(I24751), .ZN(I24752) );
NAND2_X4 U_I24753 ( .A1(g14609), .A2(I24751), .ZN(I24753) );
NAND2_X4 U_g18637 ( .A1(I24752), .A2(I24753), .ZN(g18637) );
NAND2_X4 U_I24763 ( .A1(g6194), .A2(g14573), .ZN(I24763) );
NAND2_X4 U_I24764 ( .A1(g6194), .A2(I24763), .ZN(I24764) );
NAND2_X4 U_I24765 ( .A1(g14573), .A2(I24763), .ZN(I24765) );
NAND2_X4 U_g18644 ( .A1(I24764), .A2(I24765), .ZN(g18644) );
NAND2_X4 U_g18977 ( .A1(g15797), .A2(g3006), .ZN(g18977) );
NAND2_X4 U_I25030 ( .A1(g8029), .A2(g13507), .ZN(I25030) );
NAND2_X4 U_I25031 ( .A1(g8029), .A2(I25030), .ZN(I25031) );
NAND2_X4 U_I25032 ( .A1(g13507), .A2(I25030), .ZN(I25032) );
NAND2_X4 U_g18980 ( .A1(I25031), .A2(I25032), .ZN(g18980) );
NAND2_X4 U_g19067 ( .A1(g16554), .A2(g16578), .ZN(g19067) );
NAND2_X4 U_g19084 ( .A1(g16586), .A2(g16602), .ZN(g19084) );
NAND2_X4 U_g19103 ( .A1(g18590), .A2(g2924), .ZN(g19103) );
NAND2_X4 U_g19121 ( .A1(g16682), .A2(g16697), .ZN(g19121) );
NAND2_X4 U_g19128 ( .A1(g16708), .A2(g16728), .ZN(g19128) );
NAND2_X4 U_g19135 ( .A1(g16739), .A2(g16770), .ZN(g19135) );
NAND2_X4 U_g19138 ( .A1(g16781), .A2(g16797), .ZN(g19138) );
NAND2_X4 U_g19141 ( .A1(g3088), .A2(g16825), .ZN(g19141) );
NAND2_X4 U_g19152 ( .A1(g5378), .A2(g18884), .ZN(g19152) );
NAND2_X4 U_I25532 ( .A1(g52), .A2(g18179), .ZN(I25532) );
NAND2_X4 U_I25533 ( .A1(g52), .A2(I25532), .ZN(I25533) );
NAND2_X4 U_I25534 ( .A1(g18179), .A2(I25532), .ZN(I25534) );
NAND2_X4 U_g19261 ( .A1(I25533), .A2(I25534), .ZN(g19261) );
NAND2_X4 U_I25539 ( .A1(g92), .A2(g18174), .ZN(I25539) );
NAND2_X4 U_I25540 ( .A1(g92), .A2(I25539), .ZN(I25540) );
NAND2_X4 U_I25541 ( .A1(g18174), .A2(I25539), .ZN(I25541) );
NAND2_X4 U_g19262 ( .A1(I25540), .A2(I25541), .ZN(g19262) );
NAND2_X4 U_I25560 ( .A1(g56), .A2(g17724), .ZN(I25560) );
NAND2_X4 U_I25561 ( .A1(g56), .A2(I25560), .ZN(I25561) );
NAND2_X4 U_I25562 ( .A1(g17724), .A2(I25560), .ZN(I25562) );
NAND2_X4 U_g19271 ( .A1(I25561), .A2(I25562), .ZN(g19271) );
NAND2_X4 U_I25571 ( .A1(g740), .A2(g18286), .ZN(I25571) );
NAND2_X4 U_I25572 ( .A1(g740), .A2(I25571), .ZN(I25572) );
NAND2_X4 U_I25573 ( .A1(g18286), .A2(I25571), .ZN(I25573) );
NAND2_X4 U_g19276 ( .A1(I25572), .A2(I25573), .ZN(g19276) );
NAND2_X4 U_I25578 ( .A1(g780), .A2(g18281), .ZN(I25578) );
NAND2_X4 U_I25579 ( .A1(g780), .A2(I25578), .ZN(I25579) );
NAND2_X4 U_I25580 ( .A1(g18281), .A2(I25578), .ZN(I25580) );
NAND2_X4 U_g19277 ( .A1(I25579), .A2(I25580), .ZN(g19277) );
NAND2_X4 U_I25595 ( .A1(g61), .A2(g18074), .ZN(I25595) );
NAND2_X4 U_I25596 ( .A1(g61), .A2(I25595), .ZN(I25596) );
NAND2_X4 U_I25597 ( .A1(g18074), .A2(I25595), .ZN(I25597) );
NAND2_X4 U_g19286 ( .A1(I25596), .A2(I25597), .ZN(g19286) );
NAND3_X4 U_g19288 ( .A1(g14685), .A2(g8580), .A3(g17057), .ZN(g19288) );
NAND2_X4 U_I25605 ( .A1(g744), .A2(g17825), .ZN(I25605) );
NAND2_X4 U_I25606 ( .A1(g744), .A2(I25605), .ZN(I25606) );
NAND2_X4 U_I25607 ( .A1(g17825), .A2(I25605), .ZN(I25607) );
NAND2_X4 U_g19290 ( .A1(I25606), .A2(I25607), .ZN(g19290) );
NAND2_X4 U_I25616 ( .A1(g1426), .A2(g18379), .ZN(I25616) );
NAND2_X4 U_I25617 ( .A1(g1426), .A2(I25616), .ZN(I25617) );
NAND2_X4 U_I25618 ( .A1(g18379), .A2(I25616), .ZN(I25618) );
NAND2_X4 U_g19295 ( .A1(I25617), .A2(I25618), .ZN(g19295) );
NAND2_X4 U_I25623 ( .A1(g1466), .A2(g18374), .ZN(I25623) );
NAND2_X4 U_I25624 ( .A1(g1466), .A2(I25623), .ZN(I25624) );
NAND2_X4 U_I25625 ( .A1(g18374), .A2(I25623), .ZN(I25625) );
NAND2_X4 U_g19296 ( .A1(I25624), .A2(I25625), .ZN(g19296) );
NAND2_X4 U_I25633 ( .A1(g65), .A2(g17640), .ZN(I25633) );
NAND2_X4 U_I25634 ( .A1(g65), .A2(I25633), .ZN(I25634) );
NAND2_X4 U_I25635 ( .A1(g17640), .A2(I25633), .ZN(I25635) );
NAND2_X4 U_g19300 ( .A1(I25634), .A2(I25635), .ZN(g19300) );
NAND2_X4 U_I25643 ( .A1(g749), .A2(g18190), .ZN(I25643) );
NAND2_X4 U_I25644 ( .A1(g749), .A2(I25643), .ZN(I25644) );
NAND2_X4 U_I25645 ( .A1(g18190), .A2(I25643), .ZN(I25645) );
NAND2_X4 U_g19304 ( .A1(I25644), .A2(I25645), .ZN(g19304) );
NAND3_X4 U_g19306 ( .A1(g14719), .A2(g8587), .A3(g17092), .ZN(g19306) );
NAND2_X4 U_I25653 ( .A1(g1430), .A2(g17937), .ZN(I25653) );
NAND2_X4 U_I25654 ( .A1(g1430), .A2(I25653), .ZN(I25654) );
NAND2_X4 U_I25655 ( .A1(g17937), .A2(I25653), .ZN(I25655) );
NAND2_X4 U_g19308 ( .A1(I25654), .A2(I25655), .ZN(g19308) );
NAND2_X4 U_I25664 ( .A1(g2120), .A2(g18474), .ZN(I25664) );
NAND2_X4 U_I25665 ( .A1(g2120), .A2(I25664), .ZN(I25665) );
NAND2_X4 U_I25666 ( .A1(g18474), .A2(I25664), .ZN(I25666) );
NAND2_X4 U_g19313 ( .A1(I25665), .A2(I25666), .ZN(g19313) );
NAND2_X4 U_I25671 ( .A1(g2160), .A2(g18469), .ZN(I25671) );
NAND2_X4 U_I25672 ( .A1(g2160), .A2(I25671), .ZN(I25672) );
NAND2_X4 U_I25673 ( .A1(g18469), .A2(I25671), .ZN(I25673) );
NAND2_X4 U_g19314 ( .A1(I25672), .A2(I25673), .ZN(g19314) );
NAND2_X4 U_I25681 ( .A1(g70), .A2(g17974), .ZN(I25681) );
NAND2_X4 U_I25682 ( .A1(g70), .A2(I25681), .ZN(I25682) );
NAND2_X4 U_I25683 ( .A1(g17974), .A2(I25681), .ZN(I25683) );
NAND2_X4 U_g19318 ( .A1(I25682), .A2(I25683), .ZN(g19318) );
NAND2_X4 U_I25690 ( .A1(g753), .A2(g17741), .ZN(I25690) );
NAND2_X4 U_I25691 ( .A1(g753), .A2(I25690), .ZN(I25691) );
NAND2_X4 U_I25692 ( .A1(g17741), .A2(I25690), .ZN(I25692) );
NAND2_X4 U_g19321 ( .A1(I25691), .A2(I25692), .ZN(g19321) );
NAND2_X4 U_I25700 ( .A1(g1435), .A2(g18297), .ZN(I25700) );
NAND2_X4 U_I25701 ( .A1(g1435), .A2(I25700), .ZN(I25701) );
NAND2_X4 U_I25702 ( .A1(g18297), .A2(I25700), .ZN(I25702) );
NAND2_X4 U_g19325 ( .A1(I25701), .A2(I25702), .ZN(g19325) );
NAND3_X4 U_g19327 ( .A1(g14747), .A2(g8594), .A3(g17130), .ZN(g19327) );
NAND2_X4 U_I25710 ( .A1(g2124), .A2(g18048), .ZN(I25710) );
NAND2_X4 U_I25711 ( .A1(g2124), .A2(I25710), .ZN(I25711) );
NAND2_X4 U_I25712 ( .A1(g18048), .A2(I25710), .ZN(I25712) );
NAND2_X4 U_g19329 ( .A1(I25711), .A2(I25712), .ZN(g19329) );
NAND2_X4 U_I25721 ( .A1(g74), .A2(g18341), .ZN(I25721) );
NAND2_X4 U_I25722 ( .A1(g74), .A2(I25721), .ZN(I25722) );
NAND2_X4 U_I25723 ( .A1(g18341), .A2(I25721), .ZN(I25723) );
NAND2_X4 U_g19334 ( .A1(I25722), .A2(I25723), .ZN(g19334) );
NAND2_X4 U_I25731 ( .A1(g758), .A2(g18091), .ZN(I25731) );
NAND2_X4 U_I25732 ( .A1(g758), .A2(I25731), .ZN(I25732) );
NAND2_X4 U_I25733 ( .A1(g18091), .A2(I25731), .ZN(I25733) );
NAND2_X4 U_g19345 ( .A1(I25732), .A2(I25733), .ZN(g19345) );
NAND2_X4 U_I25740 ( .A1(g1439), .A2(g17842), .ZN(I25740) );
NAND2_X4 U_I25741 ( .A1(g1439), .A2(I25740), .ZN(I25741) );
NAND2_X4 U_I25742 ( .A1(g17842), .A2(I25740), .ZN(I25742) );
NAND2_X4 U_g19348 ( .A1(I25741), .A2(I25742), .ZN(g19348) );
NAND2_X4 U_I25750 ( .A1(g2129), .A2(g18390), .ZN(I25750) );
NAND2_X4 U_I25751 ( .A1(g2129), .A2(I25750), .ZN(I25751) );
NAND2_X4 U_I25752 ( .A1(g18390), .A2(I25750), .ZN(I25752) );
NAND2_X4 U_g19352 ( .A1(I25751), .A2(I25752), .ZN(g19352) );
NAND3_X4 U_g19354 ( .A1(g14768), .A2(g8605), .A3(g17157), .ZN(g19354) );
NAND2_X4 U_I25761 ( .A1(g79), .A2(g17882), .ZN(I25761) );
NAND2_X4 U_I25762 ( .A1(g79), .A2(I25761), .ZN(I25762) );
NAND2_X4 U_I25763 ( .A1(g17882), .A2(I25761), .ZN(I25763) );
NAND2_X4 U_g19357 ( .A1(I25762), .A2(I25763), .ZN(g19357) );
NAND2_X4 U_I25771 ( .A1(g762), .A2(g18436), .ZN(I25771) );
NAND2_X4 U_I25772 ( .A1(g762), .A2(I25771), .ZN(I25772) );
NAND2_X4 U_I25773 ( .A1(g18436), .A2(I25771), .ZN(I25773) );
NAND2_X4 U_g19368 ( .A1(I25772), .A2(I25773), .ZN(g19368) );
NAND2_X4 U_I25781 ( .A1(g1444), .A2(g18207), .ZN(I25781) );
NAND2_X4 U_I25782 ( .A1(g1444), .A2(I25781), .ZN(I25782) );
NAND2_X4 U_I25783 ( .A1(g18207), .A2(I25781), .ZN(I25783) );
NAND2_X4 U_g19379 ( .A1(I25782), .A2(I25783), .ZN(g19379) );
NAND2_X4 U_I25790 ( .A1(g2133), .A2(g17954), .ZN(I25790) );
NAND2_X4 U_I25791 ( .A1(g2133), .A2(I25790), .ZN(I25791) );
NAND2_X4 U_I25792 ( .A1(g17954), .A2(I25790), .ZN(I25792) );
NAND2_X4 U_g19382 ( .A1(I25791), .A2(I25792), .ZN(g19382) );
NAND2_X4 U_I25800 ( .A1(g83), .A2(g18265), .ZN(I25800) );
NAND2_X4 U_I25801 ( .A1(g83), .A2(I25800), .ZN(I25801) );
NAND2_X4 U_I25802 ( .A1(g18265), .A2(I25800), .ZN(I25802) );
NAND2_X4 U_g19386 ( .A1(I25801), .A2(I25802), .ZN(g19386) );
NAND2_X4 U_I25809 ( .A1(g767), .A2(g17993), .ZN(I25809) );
NAND2_X4 U_I25810 ( .A1(g767), .A2(I25809), .ZN(I25810) );
NAND2_X4 U_I25811 ( .A1(g17993), .A2(I25809), .ZN(I25811) );
NAND2_X4 U_g19389 ( .A1(I25810), .A2(I25811), .ZN(g19389) );
NAND2_X4 U_I25819 ( .A1(g1448), .A2(g18509), .ZN(I25819) );
NAND2_X4 U_I25820 ( .A1(g1448), .A2(I25819), .ZN(I25820) );
NAND2_X4 U_I25821 ( .A1(g18509), .A2(I25819), .ZN(I25821) );
NAND2_X4 U_g19400 ( .A1(I25820), .A2(I25821), .ZN(g19400) );
NAND2_X4 U_I25829 ( .A1(g2138), .A2(g18314), .ZN(I25829) );
NAND2_X4 U_I25830 ( .A1(g2138), .A2(I25829), .ZN(I25830) );
NAND2_X4 U_I25831 ( .A1(g18314), .A2(I25829), .ZN(I25831) );
NAND2_X4 U_g19411 ( .A1(I25830), .A2(I25831), .ZN(g19411) );
NAND2_X4 U_I25838 ( .A1(g88), .A2(g17802), .ZN(I25838) );
NAND2_X4 U_I25839 ( .A1(g88), .A2(I25838), .ZN(I25839) );
NAND2_X4 U_I25840 ( .A1(g17802), .A2(I25838), .ZN(I25840) );
NAND2_X4 U_g19414 ( .A1(I25839), .A2(I25840), .ZN(g19414) );
NAND2_X4 U_I25846 ( .A1(g771), .A2(g18358), .ZN(I25846) );
NAND2_X4 U_I25847 ( .A1(g771), .A2(I25846), .ZN(I25847) );
NAND2_X4 U_I25848 ( .A1(g18358), .A2(I25846), .ZN(I25848) );
NAND2_X4 U_g19416 ( .A1(I25847), .A2(I25848), .ZN(g19416) );
NAND2_X4 U_I25855 ( .A1(g1453), .A2(g18110), .ZN(I25855) );
NAND2_X4 U_I25856 ( .A1(g1453), .A2(I25855), .ZN(I25856) );
NAND2_X4 U_I25857 ( .A1(g18110), .A2(I25855), .ZN(I25857) );
NAND2_X4 U_g19419 ( .A1(I25856), .A2(I25857), .ZN(g19419) );
NAND2_X4 U_I25865 ( .A1(g2142), .A2(g18573), .ZN(I25865) );
NAND2_X4 U_I25866 ( .A1(g2142), .A2(I25865), .ZN(I25866) );
NAND2_X4 U_I25867 ( .A1(g18573), .A2(I25865), .ZN(I25867) );
NAND2_X4 U_g19430 ( .A1(I25866), .A2(I25867), .ZN(g19430) );
NAND2_X4 U_I25880 ( .A1(g776), .A2(g17914), .ZN(I25880) );
NAND2_X4 U_I25881 ( .A1(g776), .A2(I25880), .ZN(I25881) );
NAND2_X4 U_I25882 ( .A1(g17914), .A2(I25880), .ZN(I25882) );
NAND2_X4 U_g19451 ( .A1(I25881), .A2(I25882), .ZN(g19451) );
NAND2_X4 U_I25888 ( .A1(g1457), .A2(g18453), .ZN(I25888) );
NAND2_X4 U_I25889 ( .A1(g1457), .A2(I25888), .ZN(I25889) );
NAND2_X4 U_I25890 ( .A1(g18453), .A2(I25888), .ZN(I25890) );
NAND2_X4 U_g19453 ( .A1(I25889), .A2(I25890), .ZN(g19453) );
NAND2_X4 U_I25897 ( .A1(g2147), .A2(g18226), .ZN(I25897) );
NAND2_X4 U_I25898 ( .A1(g2147), .A2(I25897), .ZN(I25898) );
NAND2_X4 U_I25899 ( .A1(g18226), .A2(I25897), .ZN(I25899) );
NAND2_X4 U_g19456 ( .A1(I25898), .A2(I25899), .ZN(g19456) );
NAND2_X4 U_I25913 ( .A1(g1462), .A2(g18025), .ZN(I25913) );
NAND2_X4 U_I25914 ( .A1(g1462), .A2(I25913), .ZN(I25914) );
NAND2_X4 U_I25915 ( .A1(g18025), .A2(I25913), .ZN(I25915) );
NAND2_X4 U_g19478 ( .A1(I25914), .A2(I25915), .ZN(g19478) );
NAND2_X4 U_I25921 ( .A1(g2151), .A2(g18526), .ZN(I25921) );
NAND2_X4 U_I25922 ( .A1(g2151), .A2(I25921), .ZN(I25922) );
NAND2_X4 U_I25923 ( .A1(g18526), .A2(I25921), .ZN(I25923) );
NAND2_X4 U_g19480 ( .A1(I25922), .A2(I25923), .ZN(g19480) );
NAND2_X4 U_I25938 ( .A1(g2156), .A2(g18142), .ZN(I25938) );
NAND2_X4 U_I25939 ( .A1(g2156), .A2(I25938), .ZN(I25939) );
NAND2_X4 U_I25940 ( .A1(g18142), .A2(I25938), .ZN(I25940) );
NAND2_X4 U_g19501 ( .A1(I25939), .A2(I25940), .ZN(g19501) );
NAND2_X4 U_g19865 ( .A1(g16607), .A2(g9636), .ZN(g19865) );
NAND2_X4 U_g19896 ( .A1(g16625), .A2(g9782), .ZN(g19896) );
NAND2_X4 U_g19921 ( .A1(g16639), .A2(g9928), .ZN(g19921) );
NAND2_X4 U_g19936 ( .A1(g16650), .A2(g10082), .ZN(g19936) );
NAND2_X4 U_g19954 ( .A1(g17186), .A2(g92), .ZN(g19954) );
NAND2_X4 U_g19984 ( .A1(g17197), .A2(g780), .ZN(g19984) );
NAND2_X4 U_g20022 ( .A1(g17204), .A2(g1466), .ZN(g20022) );
NAND2_X4 U_g20064 ( .A1(g17209), .A2(g2160), .ZN(g20064) );
NAND2_X4 U_g20473 ( .A1(g18085), .A2(g646), .ZN(g20473) );
NAND2_X4 U_g20481 ( .A1(g18201), .A2(g1332), .ZN(g20481) );
NAND2_X4 U_g20487 ( .A1(g18308), .A2(g2026), .ZN(g20487) );
NAND2_X4 U_g20493 ( .A1(g18401), .A2(g2720), .ZN(g20493) );
NAND2_X4 U_g20497 ( .A1(g5410), .A2(g18886), .ZN(g20497) );
NAND2_X4 U_g20522 ( .A1(g16501), .A2(g16515), .ZN(g20522) );
NAND2_X4 U_g20537 ( .A1(g18626), .A2(g3036), .ZN(g20537) );
NAND2_X4 U_g20542 ( .A1(g16523), .A2(g16546), .ZN(g20542) );
NAND2_X4 U_g20633 ( .A1(g20164), .A2(g3254), .ZN(g20633) );
NAND2_X4 U_g20648 ( .A1(g20164), .A2(g3254), .ZN(g20648) );
NAND2_X4 U_g20658 ( .A1(g20198), .A2(g3410), .ZN(g20658) );
NAND2_X4 U_g20672 ( .A1(g20164), .A2(g3254), .ZN(g20672) );
NAND2_X4 U_g20683 ( .A1(g20198), .A2(g3410), .ZN(g20683) );
NAND2_X4 U_g20693 ( .A1(g20228), .A2(g3566), .ZN(g20693) );
NAND2_X4 U_g20700 ( .A1(g20153), .A2(g2903), .ZN(g20700) );
NAND2_X4 U_g20703 ( .A1(g20164), .A2(g3254), .ZN(g20703) );
NAND2_X4 U_g20707 ( .A1(g20198), .A2(g3410), .ZN(g20707) );
NAND2_X4 U_g20718 ( .A1(g20228), .A2(g3566), .ZN(g20718) );
NAND2_X4 U_g20728 ( .A1(g20255), .A2(g3722), .ZN(g20728) );
NAND2_X4 U_g20738 ( .A1(g20198), .A2(g3410), .ZN(g20738) );
NAND2_X4 U_g20742 ( .A1(g20228), .A2(g3566), .ZN(g20742) );
NAND2_X4 U_g20753 ( .A1(g20255), .A2(g3722), .ZN(g20753) );
NAND2_X4 U_g20775 ( .A1(g20228), .A2(g3566), .ZN(g20775) );
NAND2_X4 U_g20779 ( .A1(g20255), .A2(g3722), .ZN(g20779) );
NAND2_X4 U_g20805 ( .A1(g20255), .A2(g3722), .ZN(g20805) );
NAND2_X4 U_g20825 ( .A1(g19219), .A2(g15959), .ZN(g20825) );
NAND2_X4 U_g21659 ( .A1(g20164), .A2(g6314), .ZN(g21659) );
NAND2_X4 U_I28189 ( .A1(g14079), .A2(g19444), .ZN(I28189) );
NAND2_X4 U_I28190 ( .A1(g14079), .A2(I28189), .ZN(I28190) );
NAND2_X4 U_I28191 ( .A1(g19444), .A2(I28189), .ZN(I28191) );
NAND2_X4 U_g21660 ( .A1(I28190), .A2(I28191), .ZN(g21660) );
NAND2_X4 U_g21685 ( .A1(g20164), .A2(g6232), .ZN(g21685) );
NAND2_X4 U_g21686 ( .A1(g20164), .A2(g6314), .ZN(g21686) );
NAND2_X4 U_g21688 ( .A1(g20198), .A2(g6519), .ZN(g21688) );
NAND2_X4 U_I28217 ( .A1(g14194), .A2(g19471), .ZN(I28217) );
NAND2_X4 U_I28218 ( .A1(g14194), .A2(I28217), .ZN(I28218) );
NAND2_X4 U_I28219 ( .A1(g19471), .A2(I28217), .ZN(I28219) );
NAND2_X4 U_g21689 ( .A1(I28218), .A2(I28219), .ZN(g21689) );
NAND2_X4 U_g21714 ( .A1(g20164), .A2(g6232), .ZN(g21714) );
NAND2_X4 U_g21715 ( .A1(g20164), .A2(g6314), .ZN(g21715) );
NAND4_X4 U_g21720 ( .A1(g14256), .A2(g15177), .A3(g19871), .A4(g19842), .ZN(g21720) );
NAND2_X4 U_g21721 ( .A1(g20198), .A2(g6369), .ZN(g21721) );
NAND2_X4 U_g21722 ( .A1(g20198), .A2(g6519), .ZN(g21722) );
NAND2_X4 U_g21724 ( .A1(g20228), .A2(g6783), .ZN(g21724) );
NAND2_X4 U_I28247 ( .A1(g14309), .A2(g19494), .ZN(I28247) );
NAND2_X4 U_I28248 ( .A1(g14309), .A2(I28247), .ZN(I28248) );
NAND2_X4 U_I28249 ( .A1(g19494), .A2(I28247), .ZN(I28249) );
NAND2_X4 U_g21725 ( .A1(I28248), .A2(I28249), .ZN(g21725) );
NAND2_X4 U_g21736 ( .A1(g20164), .A2(g6232), .ZN(g21736) );
NAND2_X4 U_g21737 ( .A1(g20164), .A2(g6314), .ZN(g21737) );
NAND2_X4 U_g21740 ( .A1(g20198), .A2(g6369), .ZN(g21740) );
NAND2_X4 U_g21741 ( .A1(g20198), .A2(g6519), .ZN(g21741) );
NAND4_X4 U_g21746 ( .A1(g14378), .A2(g15263), .A3(g19902), .A4(g19875), .ZN(g21746) );
NAND2_X4 U_g21747 ( .A1(g20228), .A2(g6574), .ZN(g21747) );
NAND2_X4 U_g21748 ( .A1(g20228), .A2(g6783), .ZN(g21748) );
NAND2_X4 U_g21750 ( .A1(g20255), .A2(g7085), .ZN(g21750) );
NAND2_X4 U_I28271 ( .A1(g14431), .A2(g19515), .ZN(I28271) );
NAND2_X4 U_I28272 ( .A1(g14431), .A2(I28271), .ZN(I28272) );
NAND2_X4 U_I28273 ( .A1(g19515), .A2(I28271), .ZN(I28273) );
NAND2_X4 U_g21751 ( .A1(I28272), .A2(I28273), .ZN(g21751) );
NAND2_X4 U_g21759 ( .A1(g20164), .A2(g6232), .ZN(g21759) );
NAND2_X4 U_g21760 ( .A1(g20198), .A2(g6369), .ZN(g21760) );
NAND2_X4 U_g21761 ( .A1(g20198), .A2(g6519), .ZN(g21761) );
NAND2_X4 U_g21764 ( .A1(g20228), .A2(g6574), .ZN(g21764) );
NAND2_X4 U_g21765 ( .A1(g20228), .A2(g6783), .ZN(g21765) );
NAND4_X4 U_g21770 ( .A1(g14490), .A2(g15355), .A3(g19927), .A4(g19906), .ZN(g21770) );
NAND2_X4 U_g21771 ( .A1(g20255), .A2(g6838), .ZN(g21771) );
NAND2_X4 U_g21772 ( .A1(g20255), .A2(g7085), .ZN(g21772) );
NAND2_X4 U_g21775 ( .A1(g20198), .A2(g6369), .ZN(g21775) );
NAND2_X4 U_g21776 ( .A1(g20228), .A2(g6574), .ZN(g21776) );
NAND2_X4 U_g21777 ( .A1(g20228), .A2(g6783), .ZN(g21777) );
NAND2_X4 U_g21780 ( .A1(g20255), .A2(g6838), .ZN(g21780) );
NAND2_X4 U_g21781 ( .A1(g20255), .A2(g7085), .ZN(g21781) );
NAND4_X4 U_g21786 ( .A1(g14577), .A2(g15441), .A3(g19942), .A4(g19931), .ZN(g21786) );
NAND2_X4 U_g21790 ( .A1(g20228), .A2(g6574), .ZN(g21790) );
NAND2_X4 U_g21791 ( .A1(g20255), .A2(g6838), .ZN(g21791) );
NAND2_X4 U_g21792 ( .A1(g20255), .A2(g7085), .ZN(g21792) );
NAND2_X4 U_g21804 ( .A1(g20255), .A2(g6838), .ZN(g21804) );
NAND3_X4 U_g21848 ( .A1(g17807), .A2(g19181), .A3(g19186), .ZN(g21848) );
NAND3_X4 U_g21850 ( .A1(g17979), .A2(g19187), .A3(g19191), .ZN(g21850) );
NAND3_X4 U_g21855 ( .A1(g17919), .A2(g19188), .A3(g19193), .ZN(g21855) );
NAND3_X4 U_g21857 ( .A1(g18079), .A2(g19192), .A3(g19200), .ZN(g21857) );
NAND3_X4 U_g21858 ( .A1(g18096), .A2(g19194), .A3(g19202), .ZN(g21858) );
NAND3_X4 U_g21859 ( .A1(g18030), .A2(g19195), .A3(g19204), .ZN(g21859) );
NAND3_X4 U_g21860 ( .A1(g18270), .A2(g19201), .A3(g19209), .ZN(g21860) );
NAND3_X4 U_g21862 ( .A1(g18195), .A2(g19203), .A3(g19211), .ZN(g21862) );
NAND3_X4 U_g21863 ( .A1(g18212), .A2(g19205), .A3(g19213), .ZN(g21863) );
NAND3_X4 U_g21864 ( .A1(g18147), .A2(g19206), .A3(g19215), .ZN(g21864) );
NAND3_X4 U_g21865 ( .A1(g18424), .A2(g19210), .A3(g19221), .ZN(g21865) );
NAND3_X4 U_g21866 ( .A1(g18363), .A2(g19212), .A3(g19222), .ZN(g21866) );
NAND3_X4 U_g21868 ( .A1(g18302), .A2(g19214), .A3(g19224), .ZN(g21868) );
NAND3_X4 U_g21869 ( .A1(g18319), .A2(g19216), .A3(g19226), .ZN(g21869) );
NAND3_X4 U_g21870 ( .A1(g18497), .A2(g19223), .A3(g19231), .ZN(g21870) );
NAND3_X4 U_g21871 ( .A1(g18458), .A2(g19225), .A3(g19232), .ZN(g21871) );
NAND3_X4 U_g21873 ( .A1(g18395), .A2(g19227), .A3(g19234), .ZN(g21873) );
NAND3_X4 U_g21874 ( .A1(g18561), .A2(g19233), .A3(g19244), .ZN(g21874) );
NAND3_X4 U_g21875 ( .A1(g18531), .A2(g19235), .A3(g19245), .ZN(g21875) );
NAND3_X4 U_g21877 ( .A1(g18611), .A2(g19246), .A3(g19257), .ZN(g21877) );
NAND3_X4 U_g21879 ( .A1(g18419), .A2(g19250), .A3(g19263), .ZN(g21879) );
NAND3_X4 U_g21881 ( .A1(g18492), .A2(g19264), .A3(g19278), .ZN(g21881) );
NAND3_X4 U_g21885 ( .A1(g18556), .A2(g19279), .A3(g19297), .ZN(g21885) );
NAND3_X4 U_g21888 ( .A1(g18606), .A2(g19298), .A3(g19315), .ZN(g21888) );
NAND2_X4 U_g21903 ( .A1(g20008), .A2(g3013), .ZN(g21903) );
NAND3_X4 U_g21976 ( .A1(g19242), .A2(g21120), .A3(g19275), .ZN(g21976) );
NAND3_X4 U_g21983 ( .A1(g19255), .A2(g21139), .A3(g19294), .ZN(g21983) );
NAND2_X4 U_g21989 ( .A1(g21048), .A2(g18623), .ZN(g21989) );
NAND2_X4 U_g21991 ( .A1(g21501), .A2(g21536), .ZN(g21991) );
NAND3_X4 U_g21996 ( .A1(g19268), .A2(g21159), .A3(g19312), .ZN(g21996) );
NAND2_X4 U_g22002 ( .A1(g21065), .A2(g21711), .ZN(g22002) );
NAND2_X4 U_g22005 ( .A1(g21540), .A2(g21572), .ZN(g22005) );
NAND3_X4 U_g22009 ( .A1(g19283), .A2(g21179), .A3(g19333), .ZN(g22009) );
NAND2_X4 U_g22016 ( .A1(g21576), .A2(g21605), .ZN(g22016) );
NAND2_X4 U_g22021 ( .A1(g21609), .A2(g21634), .ZN(g22021) );
NAND3_X4 U_g22050 ( .A1(g19450), .A2(g21244), .A3(g19503), .ZN(g22050) );
NAND3_X4 U_g22069 ( .A1(g19477), .A2(g21253), .A3(g19522), .ZN(g22069) );
NAND2_X4 U_g22083 ( .A1(g21774), .A2(g21787), .ZN(g22083) );
NAND3_X4 U_g22093 ( .A1(g19500), .A2(g21261), .A3(g19532), .ZN(g22093) );
NAND2_X4 U_g22108 ( .A1(g21789), .A2(g21801), .ZN(g22108) );
NAND3_X4 U_g22118 ( .A1(g19521), .A2(g21269), .A3(g19542), .ZN(g22118) );
NAND2_X4 U_g22134 ( .A1(g21803), .A2(g21809), .ZN(g22134) );
NAND2_X4 U_g22157 ( .A1(g21811), .A2(g21816), .ZN(g22157) );
NAND2_X4 U_I28726 ( .A1(g21887), .A2(g13519), .ZN(I28726) );
NAND2_X4 U_I28727 ( .A1(g21887), .A2(I28726), .ZN(I28727) );
NAND2_X4 U_I28728 ( .A1(g13519), .A2(I28726), .ZN(I28728) );
NAND2_X4 U_g22188 ( .A1(I28727), .A2(I28728), .ZN(g22188) );
NAND2_X4 U_I28741 ( .A1(g21890), .A2(g13530), .ZN(I28741) );
NAND2_X4 U_I28742 ( .A1(g21890), .A2(I28741), .ZN(I28742) );
NAND2_X4 U_I28743 ( .A1(g13530), .A2(I28741), .ZN(I28743) );
NAND2_X4 U_g22197 ( .A1(I28742), .A2(I28743), .ZN(g22197) );
NAND2_X4 U_I28753 ( .A1(g21893), .A2(g13541), .ZN(I28753) );
NAND2_X4 U_I28754 ( .A1(g21893), .A2(I28753), .ZN(I28754) );
NAND2_X4 U_I28755 ( .A1(g13541), .A2(I28753), .ZN(I28755) );
NAND2_X4 U_g22203 ( .A1(I28754), .A2(I28755), .ZN(g22203) );
NAND2_X4 U_I28765 ( .A1(g21901), .A2(g13552), .ZN(I28765) );
NAND2_X4 U_I28766 ( .A1(g21901), .A2(I28765), .ZN(I28766) );
NAND2_X4 U_I28767 ( .A1(g13552), .A2(I28765), .ZN(I28767) );
NAND2_X4 U_g22209 ( .A1(I28766), .A2(I28767), .ZN(g22209) );
NAND3_X4 U_g22317 ( .A1(g21152), .A2(g21241), .A3(g21136), .ZN(g22317) );
NAND3_X4 U_g22339 ( .A1(g14442), .A2(g21149), .A3(g10694), .ZN(g22339) );
NAND3_X4 U_g22342 ( .A1(g21172), .A2(g21249), .A3(g21156), .ZN(g22342) );
NAND3_X4 U_g22362 ( .A1(g14529), .A2(g21169), .A3(g10714), .ZN(g22362) );
NAND3_X4 U_g22365 ( .A1(g21192), .A2(g21258), .A3(g21176), .ZN(g22365) );
NAND3_X4 U_g22381 ( .A1(g21211), .A2(g14442), .A3(g10694), .ZN(g22381) );
NAND3_X4 U_g22382 ( .A1(g14584), .A2(g21189), .A3(g10735), .ZN(g22382) );
NAND3_X4 U_g22385 ( .A1(g21207), .A2(g21266), .A3(g21196), .ZN(g22385) );
NAND3_X4 U_g22396 ( .A1(g21219), .A2(g14529), .A3(g10714), .ZN(g22396) );
NAND3_X4 U_g22397 ( .A1(g14618), .A2(g21204), .A3(g10754), .ZN(g22397) );
NAND3_X4 U_g22399 ( .A1(g21230), .A2(g14584), .A3(g10735), .ZN(g22399) );
NAND3_X4 U_g22400 ( .A1(g21235), .A2(g14618), .A3(g10754), .ZN(g22400) );
NAND2_X4 U_g22608 ( .A1(g20842), .A2(g20885), .ZN(g22608) );
NAND2_X4 U_g22644 ( .A1(g20850), .A2(g20904), .ZN(g22644) );
NAND2_X4 U_g22668 ( .A1(g16075), .A2(g21271), .ZN(g22668) );
NAND2_X4 U_g22680 ( .A1(g20858), .A2(g20928), .ZN(g22680) );
NAND2_X4 U_g22708 ( .A1(g16113), .A2(g21278), .ZN(g22708) );
NAND2_X4 U_g22720 ( .A1(g20866), .A2(g20956), .ZN(g22720) );
NAND2_X4 U_g22739 ( .A1(g16164), .A2(g21285), .ZN(g22739) );
NAND2_X4 U_g22771 ( .A1(g16223), .A2(g21293), .ZN(g22771) );
NAND3_X4 U_g22809 ( .A1(g21850), .A2(g21848), .A3(g21879), .ZN(g22809) );
NAND3_X4 U_g22844 ( .A1(g21865), .A2(g21860), .A3(g21857), .ZN(g22844) );
NAND2_X4 U_g22845 ( .A1(g19441), .A2(g20885), .ZN(g22845) );
NAND2_X4 U_g22846 ( .A1(g8278), .A2(g21660), .ZN(g22846) );
NAND3_X4 U_g22850 ( .A1(g21858), .A2(g21855), .A3(g21881), .ZN(g22850) );
NAND2_X4 U_g22876 ( .A1(g21238), .A2(g83), .ZN(g22876) );
NAND3_X4 U_g22879 ( .A1(g21870), .A2(g21866), .A3(g21862), .ZN(g22879) );
NAND2_X4 U_g22880 ( .A1(g19468), .A2(g20904), .ZN(g22880) );
NAND2_X4 U_g22881 ( .A1(g8287), .A2(g21689), .ZN(g22881) );
NAND3_X4 U_g22885 ( .A1(g21863), .A2(g21859), .A3(g21885), .ZN(g22885) );
NAND2_X4 U_g22911 ( .A1(g21246), .A2(g771), .ZN(g22911) );
NAND3_X4 U_g22914 ( .A1(g21874), .A2(g21871), .A3(g21868), .ZN(g22914) );
NAND2_X4 U_g22915 ( .A1(g19491), .A2(g20928), .ZN(g22915) );
NAND2_X4 U_g22916 ( .A1(g8296), .A2(g21725), .ZN(g22916) );
NAND3_X4 U_g22920 ( .A1(g21869), .A2(g21864), .A3(g21888), .ZN(g22920) );
NAND2_X4 U_g22936 ( .A1(g21255), .A2(g1457), .ZN(g22936) );
NAND3_X4 U_g22939 ( .A1(g21877), .A2(g21875), .A3(g21873), .ZN(g22939) );
NAND2_X4 U_g22940 ( .A1(g19512), .A2(g20956), .ZN(g22940) );
NAND2_X4 U_g22941 ( .A1(g8305), .A2(g21751), .ZN(g22941) );
NAND2_X4 U_g22942 ( .A1(g21263), .A2(g2151), .ZN(g22942) );
NAND2_X4 U_g22992 ( .A1(g21636), .A2(g672), .ZN(g22992) );
NAND2_X4 U_g23003 ( .A1(g21667), .A2(g1358), .ZN(g23003) );
NAND2_X4 U_g23017 ( .A1(g21696), .A2(g2052), .ZN(g23017) );
NAND2_X4 U_g23033 ( .A1(g21732), .A2(g2746), .ZN(g23033) );
NAND2_X4 U_g23320 ( .A1(g23066), .A2(g23051), .ZN(g23320) );
NAND2_X4 U_g23325 ( .A1(g23080), .A2(g23070), .ZN(g23325) );
NAND2_X4 U_g23331 ( .A1(g22999), .A2(g22174), .ZN(g23331) );
NAND2_X4 U_g23335 ( .A1(g23096), .A2(g23083), .ZN(g23335) );
NAND2_X4 U_g23340 ( .A1(g23013), .A2(g22189), .ZN(g23340) );
NAND2_X4 U_g23344 ( .A1(g23113), .A2(g23099), .ZN(g23344) );
NAND2_X4 U_g23349 ( .A1(g23029), .A2(g22198), .ZN(g23349) );
NAND2_X4 U_g23353 ( .A1(g23046), .A2(g22204), .ZN(g23353) );
NAND2_X4 U_g23360 ( .A1(g21980), .A2(g21975), .ZN(g23360) );
NAND2_X4 U_g23364 ( .A1(g21987), .A2(g21981), .ZN(g23364) );
NAND2_X4 U_g23368 ( .A1(g23135), .A2(g22288), .ZN(g23368) );
NAND2_X4 U_g23372 ( .A1(g22000), .A2(g21988), .ZN(g23372) );
NAND2_X4 U_g23376 ( .A1(g18435), .A2(g22812), .ZN(g23376) );
NAND2_X4 U_g23377 ( .A1(g21968), .A2(g22308), .ZN(g23377) );
NAND2_X4 U_g23381 ( .A1(g22013), .A2(g22001), .ZN(g23381) );
NAND2_X4 U_g23387 ( .A1(g18508), .A2(g22852), .ZN(g23387) );
NAND2_X4 U_g23388 ( .A1(g21971), .A2(g22336), .ZN(g23388) );
NAND2_X4 U_g23394 ( .A1(g18572), .A2(g22887), .ZN(g23394) );
NAND2_X4 U_g23395 ( .A1(g21973), .A2(g22361), .ZN(g23395) );
NAND2_X4 U_g23402 ( .A1(g18622), .A2(g22922), .ZN(g23402) );
NAND3_X4 U_g23478 ( .A1(g22809), .A2(g14442), .A3(g10694), .ZN(g23478) );
NAND3_X4 U_g23486 ( .A1(g22844), .A2(g14442), .A3(g10694), .ZN(g23486) );
NAND3_X4 U_g23489 ( .A1(g22850), .A2(g14529), .A3(g10714), .ZN(g23489) );
NAND3_X4 U_g23495 ( .A1(g10694), .A2(g14442), .A3(g22316), .ZN(g23495) );
NAND3_X4 U_g23502 ( .A1(g22879), .A2(g14529), .A3(g10714), .ZN(g23502) );
NAND3_X4 U_g23505 ( .A1(g22885), .A2(g14584), .A3(g10735), .ZN(g23505) );
NAND3_X4 U_g23511 ( .A1(g10714), .A2(g14529), .A3(g22341), .ZN(g23511) );
NAND3_X4 U_g23518 ( .A1(g22914), .A2(g14584), .A3(g10735), .ZN(g23518) );
NAND3_X4 U_g23521 ( .A1(g22920), .A2(g14618), .A3(g10754), .ZN(g23521) );
NAND3_X4 U_g23526 ( .A1(g10735), .A2(g14584), .A3(g22364), .ZN(g23526) );
NAND3_X4 U_g23533 ( .A1(g22939), .A2(g14618), .A3(g10754), .ZN(g23533) );
NAND3_X4 U_g23537 ( .A1(g10754), .A2(g14618), .A3(g22384), .ZN(g23537) );
NAND2_X4 U_I30790 ( .A1(g22846), .A2(g14079), .ZN(I30790) );
NAND2_X4 U_I30791 ( .A1(g22846), .A2(I30790), .ZN(I30791) );
NAND2_X4 U_I30792 ( .A1(g14079), .A2(I30790), .ZN(I30792) );
NAND2_X4 U_g23660 ( .A1(I30791), .A2(I30792), .ZN(g23660) );
NAND2_X4 U_I30868 ( .A1(g22881), .A2(g14194), .ZN(I30868) );
NAND2_X4 U_I30869 ( .A1(g22881), .A2(I30868), .ZN(I30869) );
NAND2_X4 U_I30870 ( .A1(g14194), .A2(I30868), .ZN(I30870) );
NAND2_X4 U_g23710 ( .A1(I30869), .A2(I30870), .ZN(g23710) );
NAND2_X4 U_I30952 ( .A1(g22916), .A2(g14309), .ZN(I30952) );
NAND2_X4 U_I30953 ( .A1(g22916), .A2(I30952), .ZN(I30953) );
NAND2_X4 U_I30954 ( .A1(g14309), .A2(I30952), .ZN(I30954) );
NAND2_X4 U_g23764 ( .A1(I30953), .A2(I30954), .ZN(g23764) );
NAND2_X4 U_I31035 ( .A1(g22941), .A2(g14431), .ZN(I31035) );
NAND2_X4 U_I31036 ( .A1(g22941), .A2(I31035), .ZN(I31036) );
NAND2_X4 U_I31037 ( .A1(g14431), .A2(I31035), .ZN(I31037) );
NAND2_X4 U_g23819 ( .A1(I31036), .A2(I31037), .ZN(g23819) );
NAND2_X4 U_g23906 ( .A1(g22812), .A2(g13958), .ZN(g23906) );
NAND2_X4 U_g23936 ( .A1(g22812), .A2(g13922), .ZN(g23936) );
NAND2_X4 U_g23937 ( .A1(g22812), .A2(g13918), .ZN(g23937) );
NAND2_X4 U_g23938 ( .A1(g22852), .A2(g14028), .ZN(g23938) );
NAND2_X4 U_g23953 ( .A1(g22812), .A2(g14525), .ZN(g23953) );
NAND2_X4 U_g23968 ( .A1(g22852), .A2(g13978), .ZN(g23968) );
NAND2_X4 U_g23969 ( .A1(g22852), .A2(g13974), .ZN(g23969) );
NAND2_X4 U_g23970 ( .A1(g22887), .A2(g14119), .ZN(g23970) );
NAND2_X4 U_g23973 ( .A1(g22812), .A2(g14450), .ZN(g23973) );
NAND2_X4 U_g23982 ( .A1(g22852), .A2(g14580), .ZN(g23982) );
NAND2_X4 U_g23997 ( .A1(g22887), .A2(g14048), .ZN(g23997) );
NAND2_X4 U_g23998 ( .A1(g22887), .A2(g14044), .ZN(g23998) );
NAND2_X4 U_g23999 ( .A1(g22922), .A2(g14234), .ZN(g23999) );
NAND2_X4 U_g24002 ( .A1(g22812), .A2(g14355), .ZN(g24002) );
NAND2_X4 U_g24003 ( .A1(g22852), .A2(g14537), .ZN(g24003) );
NAND2_X4 U_g24012 ( .A1(g22887), .A2(g14614), .ZN(g24012) );
NAND2_X4 U_g24027 ( .A1(g22922), .A2(g14139), .ZN(g24027) );
NAND2_X4 U_g24028 ( .A1(g22922), .A2(g14135), .ZN(g24028) );
NAND2_X4 U_g24034 ( .A1(g22812), .A2(g14252), .ZN(g24034) );
NAND2_X4 U_g24036 ( .A1(g22852), .A2(g14467), .ZN(g24036) );
NAND2_X4 U_g24037 ( .A1(g22887), .A2(g14592), .ZN(g24037) );
NAND2_X4 U_g24046 ( .A1(g22922), .A2(g14637), .ZN(g24046) );
NAND2_X4 U_g24052 ( .A1(g22812), .A2(g14171), .ZN(g24052) );
NAND2_X4 U_g24054 ( .A1(g22852), .A2(g14374), .ZN(g24054) );
NAND2_X4 U_g24056 ( .A1(g22887), .A2(g14554), .ZN(g24056) );
NAND2_X4 U_g24057 ( .A1(g22922), .A2(g14626), .ZN(g24057) );
NAND2_X4 U_g24058 ( .A1(g22812), .A2(g14086), .ZN(g24058) );
NAND2_X4 U_g24065 ( .A1(g22852), .A2(g14286), .ZN(g24065) );
NAND2_X4 U_g24067 ( .A1(g22887), .A2(g14486), .ZN(g24067) );
NAND2_X4 U_g24069 ( .A1(g22922), .A2(g14609), .ZN(g24069) );
NAND2_X4 U_g24070 ( .A1(g22812), .A2(g14011), .ZN(g24070) );
NAND2_X4 U_g24071 ( .A1(g22852), .A2(g14201), .ZN(g24071) );
NAND2_X4 U_g24078 ( .A1(g22887), .A2(g14408), .ZN(g24078) );
NAND2_X4 U_g24080 ( .A1(g22922), .A2(g14573), .ZN(g24080) );
NAND2_X4 U_g24081 ( .A1(g22852), .A2(g14102), .ZN(g24081) );
NAND2_X4 U_g24082 ( .A1(g22887), .A2(g14316), .ZN(g24082) );
NAND2_X4 U_g24089 ( .A1(g22922), .A2(g14520), .ZN(g24089) );
NAND2_X4 U_g24090 ( .A1(g22887), .A2(g14217), .ZN(g24090) );
NAND2_X4 U_g24091 ( .A1(g22922), .A2(g14438), .ZN(g24091) );
NAND2_X4 U_g24093 ( .A1(g22922), .A2(g14332), .ZN(g24093) );
NAND2_X4 U_g24100 ( .A1(g20885), .A2(g22175), .ZN(g24100) );
NAND2_X4 U_g24109 ( .A1(g20904), .A2(g22190), .ZN(g24109) );
NAND2_X4 U_g24126 ( .A1(g20928), .A2(g22199), .ZN(g24126) );
NAND2_X4 U_g24145 ( .A1(g20956), .A2(g22205), .ZN(g24145) );
NAND2_X4 U_g24442 ( .A1(g23644), .A2(g3306), .ZN(g24442) );
NAND2_X4 U_g24443 ( .A1(g23644), .A2(g3306), .ZN(g24443) );
NAND2_X4 U_g24444 ( .A1(g23694), .A2(g3462), .ZN(g24444) );
NAND2_X4 U_g24447 ( .A1(g23644), .A2(g3306), .ZN(g24447) );
NAND2_X4 U_g24448 ( .A1(g23923), .A2(g3338), .ZN(g24448) );
NAND2_X4 U_g24449 ( .A1(g23694), .A2(g3462), .ZN(g24449) );
NAND2_X4 U_g24450 ( .A1(g23748), .A2(g3618), .ZN(g24450) );
NAND2_X4 U_g24451 ( .A1(g23644), .A2(g3306), .ZN(g24451) );
NAND2_X4 U_g24452 ( .A1(g23923), .A2(g3338), .ZN(g24452) );
NAND2_X4 U_g24453 ( .A1(g23694), .A2(g3462), .ZN(g24453) );
NAND2_X4 U_g24454 ( .A1(g23955), .A2(g3494), .ZN(g24454) );
NAND2_X4 U_g24455 ( .A1(g23748), .A2(g3618), .ZN(g24455) );
NAND2_X4 U_g24456 ( .A1(g23803), .A2(g3774), .ZN(g24456) );
NAND2_X4 U_g24457 ( .A1(g23923), .A2(g3338), .ZN(g24457) );
NAND2_X4 U_g24458 ( .A1(g23694), .A2(g3462), .ZN(g24458) );
NAND2_X4 U_g24459 ( .A1(g23955), .A2(g3494), .ZN(g24459) );
NAND2_X4 U_g24460 ( .A1(g23748), .A2(g3618), .ZN(g24460) );
NAND2_X4 U_g24461 ( .A1(g23984), .A2(g3650), .ZN(g24461) );
NAND2_X4 U_g24462 ( .A1(g23803), .A2(g3774), .ZN(g24462) );
NAND2_X4 U_g24463 ( .A1(g23923), .A2(g3338), .ZN(g24463) );
NAND2_X4 U_g24464 ( .A1(g23955), .A2(g3494), .ZN(g24464) );
NAND2_X4 U_g24465 ( .A1(g23748), .A2(g3618), .ZN(g24465) );
NAND2_X4 U_g24466 ( .A1(g23984), .A2(g3650), .ZN(g24466) );
NAND2_X4 U_g24467 ( .A1(g23803), .A2(g3774), .ZN(g24467) );
NAND2_X4 U_g24468 ( .A1(g24014), .A2(g3806), .ZN(g24468) );
NAND2_X4 U_g24469 ( .A1(g23955), .A2(g3494), .ZN(g24469) );
NAND2_X4 U_g24470 ( .A1(g23984), .A2(g3650), .ZN(g24470) );
NAND2_X4 U_g24471 ( .A1(g23803), .A2(g3774), .ZN(g24471) );
NAND2_X4 U_g24472 ( .A1(g24014), .A2(g3806), .ZN(g24472) );
NAND2_X4 U_g24474 ( .A1(g23984), .A2(g3650), .ZN(g24474) );
NAND2_X4 U_g24475 ( .A1(g24014), .A2(g3806), .ZN(g24475) );
NAND2_X4 U_g24477 ( .A1(g24014), .A2(g3806), .ZN(g24477) );
NAND2_X4 U_g24616 ( .A1(g499), .A2(g23376), .ZN(g24616) );
NAND2_X4 U_g24627 ( .A1(g1186), .A2(g23387), .ZN(g24627) );
NAND2_X4 U_g24641 ( .A1(g1880), .A2(g23394), .ZN(g24641) );
NAND2_X4 U_g24660 ( .A1(g2574), .A2(g23402), .ZN(g24660) );
NAND2_X4 U_I32265 ( .A1(g17903), .A2(g23936), .ZN(I32265) );
NAND2_X4 U_I32266 ( .A1(g17903), .A2(I32265), .ZN(I32266) );
NAND2_X4 U_I32267 ( .A1(g23936), .A2(I32265), .ZN(I32267) );
NAND2_X4 U_g24753 ( .A1(I32266), .A2(I32267), .ZN(g24753) );
NAND2_X4 U_I32284 ( .A1(g17815), .A2(g23953), .ZN(I32284) );
NAND2_X4 U_I32285 ( .A1(g17815), .A2(I32284), .ZN(I32285) );
NAND2_X4 U_I32286 ( .A1(g23953), .A2(I32284), .ZN(I32286) );
NAND2_X4 U_g24766 ( .A1(I32285), .A2(I32286), .ZN(g24766) );
NAND2_X4 U_I32295 ( .A1(g18014), .A2(g23968), .ZN(I32295) );
NAND2_X4 U_I32296 ( .A1(g18014), .A2(I32295), .ZN(I32296) );
NAND2_X4 U_I32297 ( .A1(g23968), .A2(I32295), .ZN(I32297) );
NAND2_X4 U_g24771 ( .A1(I32296), .A2(I32297), .ZN(g24771) );
NAND2_X4 U_I32308 ( .A1(g17903), .A2(g23973), .ZN(I32308) );
NAND2_X4 U_I32309 ( .A1(g17903), .A2(I32308), .ZN(I32309) );
NAND2_X4 U_I32310 ( .A1(g23973), .A2(I32308), .ZN(I32310) );
NAND2_X4 U_g24778 ( .A1(I32309), .A2(I32310), .ZN(g24778) );
NAND2_X4 U_I32323 ( .A1(g17927), .A2(g23982), .ZN(I32323) );
NAND2_X4 U_I32324 ( .A1(g17927), .A2(I32323), .ZN(I32324) );
NAND2_X4 U_I32325 ( .A1(g23982), .A2(I32323), .ZN(I32325) );
NAND2_X4 U_g24787 ( .A1(I32324), .A2(I32325), .ZN(g24787) );
NAND2_X4 U_I32333 ( .A1(g18131), .A2(g23997), .ZN(I32333) );
NAND2_X4 U_I32334 ( .A1(g18131), .A2(I32333), .ZN(I32334) );
NAND2_X4 U_I32335 ( .A1(g23997), .A2(I32333), .ZN(I32335) );
NAND2_X4 U_g24791 ( .A1(I32334), .A2(I32335), .ZN(g24791) );
NAND2_X4 U_I32345 ( .A1(g17815), .A2(g24002), .ZN(I32345) );
NAND2_X4 U_I32346 ( .A1(g17815), .A2(I32345), .ZN(I32346) );
NAND2_X4 U_I32347 ( .A1(g24002), .A2(I32345), .ZN(I32347) );
NAND2_X4 U_g24797 ( .A1(I32346), .A2(I32347), .ZN(g24797) );
NAND2_X4 U_I32355 ( .A1(g18014), .A2(g24003), .ZN(I32355) );
NAND2_X4 U_I32356 ( .A1(g18014), .A2(I32355), .ZN(I32356) );
NAND2_X4 U_I32357 ( .A1(g24003), .A2(I32355), .ZN(I32357) );
NAND2_X4 U_g24801 ( .A1(I32356), .A2(I32357), .ZN(g24801) );
NAND2_X4 U_I32368 ( .A1(g18038), .A2(g24012), .ZN(I32368) );
NAND2_X4 U_I32369 ( .A1(g18038), .A2(I32368), .ZN(I32369) );
NAND2_X4 U_I32370 ( .A1(g24012), .A2(I32368), .ZN(I32370) );
NAND2_X4 U_g24808 ( .A1(I32369), .A2(I32370), .ZN(g24808) );
NAND2_X4 U_I32378 ( .A1(g18247), .A2(g24027), .ZN(I32378) );
NAND2_X4 U_I32379 ( .A1(g18247), .A2(I32378), .ZN(I32379) );
NAND2_X4 U_I32380 ( .A1(g24027), .A2(I32378), .ZN(I32380) );
NAND2_X4 U_g24812 ( .A1(I32379), .A2(I32380), .ZN(g24812) );
NAND2_X4 U_g24814 ( .A1(g24239), .A2(g24244), .ZN(g24814) );
NAND2_X4 U_I32391 ( .A1(g17903), .A2(g24034), .ZN(I32391) );
NAND2_X4 U_I32392 ( .A1(g17903), .A2(I32391), .ZN(I32392) );
NAND2_X4 U_I32393 ( .A1(g24034), .A2(I32391), .ZN(I32393) );
NAND2_X4 U_g24817 ( .A1(I32392), .A2(I32393), .ZN(g24817) );
NAND2_X4 U_I32400 ( .A1(g17927), .A2(g24036), .ZN(I32400) );
NAND2_X4 U_I32401 ( .A1(g17927), .A2(I32400), .ZN(I32401) );
NAND2_X4 U_I32402 ( .A1(g24036), .A2(I32400), .ZN(I32402) );
NAND2_X4 U_g24820 ( .A1(I32401), .A2(I32402), .ZN(g24820) );
NAND2_X4 U_I32409 ( .A1(g18131), .A2(g24037), .ZN(I32409) );
NAND2_X4 U_I32410 ( .A1(g18131), .A2(I32409), .ZN(I32410) );
NAND2_X4 U_I32411 ( .A1(g24037), .A2(I32409), .ZN(I32411) );
NAND2_X4 U_g24823 ( .A1(I32410), .A2(I32411), .ZN(g24823) );
NAND2_X4 U_I32422 ( .A1(g18155), .A2(g24046), .ZN(I32422) );
NAND2_X4 U_I32423 ( .A1(g18155), .A2(I32422), .ZN(I32423) );
NAND2_X4 U_I32424 ( .A1(g24046), .A2(I32422), .ZN(I32424) );
NAND2_X4 U_g24830 ( .A1(I32423), .A2(I32424), .ZN(g24830) );
NAND2_X4 U_I32430 ( .A1(g17815), .A2(g24052), .ZN(I32430) );
NAND2_X4 U_I32431 ( .A1(g17815), .A2(I32430), .ZN(I32431) );
NAND2_X4 U_I32432 ( .A1(g24052), .A2(I32430), .ZN(I32432) );
NAND2_X4 U_g24832 ( .A1(I32431), .A2(I32432), .ZN(g24832) );
NAND2_X4 U_g24833 ( .A1(g24245), .A2(g24252), .ZN(g24833) );
NAND2_X4 U_I32443 ( .A1(g18014), .A2(g24054), .ZN(I32443) );
NAND2_X4 U_I32444 ( .A1(g18014), .A2(I32443), .ZN(I32444) );
NAND2_X4 U_I32445 ( .A1(g24054), .A2(I32443), .ZN(I32445) );
NAND2_X4 U_g24837 ( .A1(I32444), .A2(I32445), .ZN(g24837) );
NAND2_X4 U_I32451 ( .A1(g18038), .A2(g24056), .ZN(I32451) );
NAND2_X4 U_I32452 ( .A1(g18038), .A2(I32451), .ZN(I32452) );
NAND2_X4 U_I32453 ( .A1(g24056), .A2(I32451), .ZN(I32453) );
NAND2_X4 U_g24839 ( .A1(I32452), .A2(I32453), .ZN(g24839) );
NAND2_X4 U_I32460 ( .A1(g18247), .A2(g24057), .ZN(I32460) );
NAND2_X4 U_I32461 ( .A1(g18247), .A2(I32460), .ZN(I32461) );
NAND2_X4 U_I32462 ( .A1(g24057), .A2(I32460), .ZN(I32462) );
NAND2_X4 U_g24842 ( .A1(I32461), .A2(I32462), .ZN(g24842) );
NAND2_X4 U_I32468 ( .A1(g17903), .A2(g24058), .ZN(I32468) );
NAND2_X4 U_I32469 ( .A1(g17903), .A2(I32468), .ZN(I32469) );
NAND2_X4 U_I32470 ( .A1(g24058), .A2(I32468), .ZN(I32470) );
NAND2_X4 U_g24844 ( .A1(I32469), .A2(I32470), .ZN(g24844) );
NAND2_X4 U_I32478 ( .A1(g17927), .A2(g24065), .ZN(I32478) );
NAND2_X4 U_I32479 ( .A1(g17927), .A2(I32478), .ZN(I32479) );
NAND2_X4 U_I32480 ( .A1(g24065), .A2(I32478), .ZN(I32480) );
NAND2_X4 U_g24848 ( .A1(I32479), .A2(I32480), .ZN(g24848) );
NAND2_X4 U_g24849 ( .A1(g24254), .A2(g24257), .ZN(g24849) );
NAND2_X4 U_I32490 ( .A1(g18131), .A2(g24067), .ZN(I32490) );
NAND2_X4 U_I32491 ( .A1(g18131), .A2(I32490), .ZN(I32491) );
NAND2_X4 U_I32492 ( .A1(g24067), .A2(I32490), .ZN(I32492) );
NAND2_X4 U_g24852 ( .A1(I32491), .A2(I32492), .ZN(g24852) );
NAND2_X4 U_I32498 ( .A1(g18155), .A2(g24069), .ZN(I32498) );
NAND2_X4 U_I32499 ( .A1(g18155), .A2(I32498), .ZN(I32499) );
NAND2_X4 U_I32500 ( .A1(g24069), .A2(I32498), .ZN(I32500) );
NAND2_X4 U_g24854 ( .A1(I32499), .A2(I32500), .ZN(g24854) );
NAND2_X4 U_I32509 ( .A1(g17815), .A2(g24070), .ZN(I32509) );
NAND2_X4 U_I32510 ( .A1(g17815), .A2(I32509), .ZN(I32510) );
NAND2_X4 U_I32511 ( .A1(g24070), .A2(I32509), .ZN(I32511) );
NAND2_X4 U_g24857 ( .A1(I32510), .A2(I32511), .ZN(g24857) );
NAND2_X4 U_I32518 ( .A1(g18014), .A2(g24071), .ZN(I32518) );
NAND2_X4 U_I32519 ( .A1(g18014), .A2(I32518), .ZN(I32519) );
NAND2_X4 U_I32520 ( .A1(g24071), .A2(I32518), .ZN(I32520) );
NAND2_X4 U_g24860 ( .A1(I32519), .A2(I32520), .ZN(g24860) );
NAND2_X4 U_I32526 ( .A1(g18038), .A2(g24078), .ZN(I32526) );
NAND2_X4 U_I32527 ( .A1(g18038), .A2(I32526), .ZN(I32527) );
NAND2_X4 U_I32528 ( .A1(g24078), .A2(I32526), .ZN(I32528) );
NAND2_X4 U_g24862 ( .A1(I32527), .A2(I32528), .ZN(g24862) );
NAND2_X4 U_g24863 ( .A1(g24258), .A2(g23319), .ZN(g24863) );
NAND2_X4 U_I32538 ( .A1(g18247), .A2(g24080), .ZN(I32538) );
NAND2_X4 U_I32539 ( .A1(g18247), .A2(I32538), .ZN(I32539) );
NAND2_X4 U_I32540 ( .A1(g24080), .A2(I32538), .ZN(I32540) );
NAND2_X4 U_g24866 ( .A1(I32539), .A2(I32540), .ZN(g24866) );
NAND2_X4 U_I32546 ( .A1(g17903), .A2(g23906), .ZN(I32546) );
NAND2_X4 U_I32547 ( .A1(g17903), .A2(I32546), .ZN(I32547) );
NAND2_X4 U_I32548 ( .A1(g23906), .A2(I32546), .ZN(I32548) );
NAND2_X4 U_g24868 ( .A1(I32547), .A2(I32548), .ZN(g24868) );
NAND2_X4 U_I32559 ( .A1(g17927), .A2(g24081), .ZN(I32559) );
NAND2_X4 U_I32560 ( .A1(g17927), .A2(I32559), .ZN(I32560) );
NAND2_X4 U_I32561 ( .A1(g24081), .A2(I32559), .ZN(I32561) );
NAND2_X4 U_g24873 ( .A1(I32560), .A2(I32561), .ZN(g24873) );
NAND2_X4 U_I32567 ( .A1(g18131), .A2(g24082), .ZN(I32567) );
NAND2_X4 U_I32568 ( .A1(g18131), .A2(I32567), .ZN(I32568) );
NAND2_X4 U_I32569 ( .A1(g24082), .A2(I32567), .ZN(I32569) );
NAND2_X4 U_g24875 ( .A1(I32568), .A2(I32569), .ZN(g24875) );
NAND2_X4 U_I32575 ( .A1(g18155), .A2(g24089), .ZN(I32575) );
NAND2_X4 U_I32576 ( .A1(g18155), .A2(I32575), .ZN(I32576) );
NAND2_X4 U_I32577 ( .A1(g24089), .A2(I32575), .ZN(I32577) );
NAND2_X4 U_g24877 ( .A1(I32576), .A2(I32577), .ZN(g24877) );
NAND2_X4 U_I32586 ( .A1(g17815), .A2(g23937), .ZN(I32586) );
NAND2_X4 U_I32587 ( .A1(g17815), .A2(I32586), .ZN(I32587) );
NAND2_X4 U_I32588 ( .A1(g23937), .A2(I32586), .ZN(I32588) );
NAND2_X4 U_g24880 ( .A1(I32587), .A2(I32588), .ZN(g24880) );
NAND2_X4 U_I32595 ( .A1(g18014), .A2(g23938), .ZN(I32595) );
NAND2_X4 U_I32596 ( .A1(g18014), .A2(I32595), .ZN(I32596) );
NAND2_X4 U_I32597 ( .A1(g23938), .A2(I32595), .ZN(I32597) );
NAND2_X4 U_g24883 ( .A1(I32596), .A2(I32597), .ZN(g24883) );
NAND2_X4 U_I32607 ( .A1(g18038), .A2(g24090), .ZN(I32607) );
NAND2_X4 U_I32608 ( .A1(g18038), .A2(I32607), .ZN(I32608) );
NAND2_X4 U_I32609 ( .A1(g24090), .A2(I32607), .ZN(I32609) );
NAND2_X4 U_g24887 ( .A1(I32608), .A2(I32609), .ZN(g24887) );
NAND2_X4 U_I32615 ( .A1(g18247), .A2(g24091), .ZN(I32615) );
NAND2_X4 U_I32616 ( .A1(g18247), .A2(I32615), .ZN(I32616) );
NAND2_X4 U_I32617 ( .A1(g24091), .A2(I32615), .ZN(I32617) );
NAND2_X4 U_g24889 ( .A1(I32616), .A2(I32617), .ZN(g24889) );
NAND2_X4 U_I32624 ( .A1(g17927), .A2(g23969), .ZN(I32624) );
NAND2_X4 U_I32625 ( .A1(g17927), .A2(I32624), .ZN(I32625) );
NAND2_X4 U_I32626 ( .A1(g23969), .A2(I32624), .ZN(I32626) );
NAND2_X4 U_g24897 ( .A1(I32625), .A2(I32626), .ZN(g24897) );
NAND2_X4 U_I32633 ( .A1(g18131), .A2(g23970), .ZN(I32633) );
NAND2_X4 U_I32634 ( .A1(g18131), .A2(I32633), .ZN(I32634) );
NAND2_X4 U_I32635 ( .A1(g23970), .A2(I32633), .ZN(I32635) );
NAND2_X4 U_g24900 ( .A1(I32634), .A2(I32635), .ZN(g24900) );
NAND2_X4 U_I32645 ( .A1(g18155), .A2(g24093), .ZN(I32645) );
NAND2_X4 U_I32646 ( .A1(g18155), .A2(I32645), .ZN(I32646) );
NAND2_X4 U_I32647 ( .A1(g24093), .A2(I32645), .ZN(I32647) );
NAND2_X4 U_g24904 ( .A1(I32646), .A2(I32647), .ZN(g24904) );
NAND2_X4 U_I32659 ( .A1(g18038), .A2(g23998), .ZN(I32659) );
NAND2_X4 U_I32660 ( .A1(g18038), .A2(I32659), .ZN(I32660) );
NAND2_X4 U_I32661 ( .A1(g23998), .A2(I32659), .ZN(I32661) );
NAND2_X4 U_g24920 ( .A1(I32660), .A2(I32661), .ZN(g24920) );
NAND2_X4 U_I32668 ( .A1(g18247), .A2(g23999), .ZN(I32668) );
NAND2_X4 U_I32669 ( .A1(g18247), .A2(I32668), .ZN(I32669) );
NAND2_X4 U_I32670 ( .A1(g23999), .A2(I32668), .ZN(I32670) );
NAND2_X4 U_g24923 ( .A1(I32669), .A2(I32670), .ZN(g24923) );
NAND2_X4 U_I32677 ( .A1(g23823), .A2(g14165), .ZN(I32677) );
NAND2_X4 U_I32678 ( .A1(g23823), .A2(I32677), .ZN(I32678) );
NAND2_X4 U_I32679 ( .A1(g14165), .A2(I32677), .ZN(I32679) );
NAND2_X4 U_g24928 ( .A1(I32678), .A2(I32679), .ZN(g24928) );
NAND2_X4 U_I32686 ( .A1(g18155), .A2(g24028), .ZN(I32686) );
NAND2_X4 U_I32687 ( .A1(g18155), .A2(I32686), .ZN(I32687) );
NAND2_X4 U_I32688 ( .A1(g24028), .A2(I32686), .ZN(I32688) );
NAND2_X4 U_g24937 ( .A1(I32687), .A2(I32688), .ZN(g24937) );
NAND2_X4 U_I32695 ( .A1(g23858), .A2(g14280), .ZN(I32695) );
NAND2_X4 U_I32696 ( .A1(g23858), .A2(I32695), .ZN(I32696) );
NAND2_X4 U_I32697 ( .A1(g14280), .A2(I32695), .ZN(I32697) );
NAND2_X4 U_g24940 ( .A1(I32696), .A2(I32697), .ZN(g24940) );
NAND2_X4 U_I32708 ( .A1(g23892), .A2(g14402), .ZN(I32708) );
NAND2_X4 U_I32709 ( .A1(g23892), .A2(I32708), .ZN(I32709) );
NAND2_X4 U_I32710 ( .A1(g14402), .A2(I32708), .ZN(I32710) );
NAND2_X4 U_g24951 ( .A1(I32709), .A2(I32710), .ZN(g24951) );
NAND2_X4 U_I32724 ( .A1(g23913), .A2(g14514), .ZN(I32724) );
NAND2_X4 U_I32725 ( .A1(g23913), .A2(I32724), .ZN(I32725) );
NAND2_X4 U_I32726 ( .A1(g14514), .A2(I32724), .ZN(I32726) );
NAND2_X4 U_g24963 ( .A1(I32725), .A2(I32726), .ZN(g24963) );
NAND2_X4 U_g24975 ( .A1(g23497), .A2(g74), .ZN(g24975) );
NAND2_X4 U_g24986 ( .A1(g23513), .A2(g762), .ZN(g24986) );
NAND2_X4 U_g24997 ( .A1(g23528), .A2(g1448), .ZN(g24997) );
NAND2_X4 U_g25004 ( .A1(g23644), .A2(g6448), .ZN(g25004) );
NAND2_X4 U_g25005 ( .A1(g23539), .A2(g2142), .ZN(g25005) );
NAND2_X4 U_g25008 ( .A1(g23644), .A2(g5438), .ZN(g25008) );
NAND2_X4 U_g25009 ( .A1(g23644), .A2(g6448), .ZN(g25009) );
NAND2_X4 U_g25010 ( .A1(g23694), .A2(g6713), .ZN(g25010) );
NAND2_X4 U_g25011 ( .A1(g23644), .A2(g5438), .ZN(g25011) );
NAND2_X4 U_g25012 ( .A1(g23644), .A2(g6448), .ZN(g25012) );
NAND2_X4 U_g25013 ( .A1(g23923), .A2(g6643), .ZN(g25013) );
NAND2_X4 U_g25014 ( .A1(g23694), .A2(g5473), .ZN(g25014) );
NAND2_X4 U_g25015 ( .A1(g23694), .A2(g6713), .ZN(g25015) );
NAND2_X4 U_g25016 ( .A1(g23748), .A2(g7015), .ZN(g25016) );
NAND2_X4 U_g25017 ( .A1(g23644), .A2(g5438), .ZN(g25017) );
NAND2_X4 U_g25018 ( .A1(g23644), .A2(g6448), .ZN(g25018) );
NAND2_X4 U_g25019 ( .A1(g23923), .A2(g6486), .ZN(g25019) );
NAND2_X4 U_g25020 ( .A1(g23923), .A2(g6643), .ZN(g25020) );
NAND2_X4 U_g25021 ( .A1(g23694), .A2(g5473), .ZN(g25021) );
NAND2_X4 U_g25022 ( .A1(g23694), .A2(g6713), .ZN(g25022) );
NAND2_X4 U_g25023 ( .A1(g23955), .A2(g6945), .ZN(g25023) );
NAND2_X4 U_g25024 ( .A1(g23748), .A2(g5512), .ZN(g25024) );
NAND2_X4 U_g25025 ( .A1(g23748), .A2(g7015), .ZN(g25025) );
NAND2_X4 U_g25026 ( .A1(g23803), .A2(g7265), .ZN(g25026) );
NAND2_X4 U_g25028 ( .A1(g23644), .A2(g5438), .ZN(g25028) );
NAND2_X4 U_g25029 ( .A1(g23923), .A2(g6486), .ZN(g25029) );
NAND2_X4 U_g25030 ( .A1(g23923), .A2(g6643), .ZN(g25030) );
NAND2_X4 U_g25031 ( .A1(g23694), .A2(g5473), .ZN(g25031) );
NAND2_X4 U_g25032 ( .A1(g23694), .A2(g6713), .ZN(g25032) );
NAND2_X4 U_g25033 ( .A1(g23955), .A2(g6751), .ZN(g25033) );
NAND2_X4 U_g25034 ( .A1(g23955), .A2(g6945), .ZN(g25034) );
NAND2_X4 U_g25035 ( .A1(g23748), .A2(g5512), .ZN(g25035) );
NAND2_X4 U_g25036 ( .A1(g23748), .A2(g7015), .ZN(g25036) );
NAND2_X4 U_g25037 ( .A1(g23984), .A2(g7195), .ZN(g25037) );
NAND2_X4 U_g25038 ( .A1(g23803), .A2(g5556), .ZN(g25038) );
NAND2_X4 U_g25039 ( .A1(g23803), .A2(g7265), .ZN(g25039) );
NAND2_X4 U_g25040 ( .A1(g23923), .A2(g6486), .ZN(g25040) );
NAND2_X4 U_g25041 ( .A1(g23923), .A2(g6643), .ZN(g25041) );
NAND2_X4 U_g25043 ( .A1(g23694), .A2(g5473), .ZN(g25043) );
NAND2_X4 U_g25044 ( .A1(g23955), .A2(g6751), .ZN(g25044) );
NAND2_X4 U_g25045 ( .A1(g23955), .A2(g6945), .ZN(g25045) );
NAND2_X4 U_g25046 ( .A1(g23748), .A2(g5512), .ZN(g25046) );
NAND2_X4 U_g25047 ( .A1(g23748), .A2(g7015), .ZN(g25047) );
NAND2_X4 U_g25048 ( .A1(g23984), .A2(g7053), .ZN(g25048) );
NAND2_X4 U_g25049 ( .A1(g23984), .A2(g7195), .ZN(g25049) );
NAND2_X4 U_g25050 ( .A1(g23803), .A2(g5556), .ZN(g25050) );
NAND2_X4 U_g25051 ( .A1(g23803), .A2(g7265), .ZN(g25051) );
NAND2_X4 U_g25052 ( .A1(g24014), .A2(g7391), .ZN(g25052) );
NAND2_X4 U_g25053 ( .A1(g23923), .A2(g6486), .ZN(g25053) );
NAND2_X4 U_g25054 ( .A1(g23955), .A2(g6751), .ZN(g25054) );
NAND2_X4 U_g25055 ( .A1(g23955), .A2(g6945), .ZN(g25055) );
NAND2_X4 U_g25057 ( .A1(g23748), .A2(g5512), .ZN(g25057) );
NAND2_X4 U_g25058 ( .A1(g23984), .A2(g7053), .ZN(g25058) );
NAND2_X4 U_g25059 ( .A1(g23984), .A2(g7195), .ZN(g25059) );
NAND2_X4 U_g25060 ( .A1(g23803), .A2(g5556), .ZN(g25060) );
NAND2_X4 U_g25061 ( .A1(g23803), .A2(g7265), .ZN(g25061) );
NAND2_X4 U_g25062 ( .A1(g24014), .A2(g7303), .ZN(g25062) );
NAND2_X4 U_g25063 ( .A1(g24014), .A2(g7391), .ZN(g25063) );
NAND2_X4 U_g25064 ( .A1(g23955), .A2(g6751), .ZN(g25064) );
NAND2_X4 U_g25065 ( .A1(g23984), .A2(g7053), .ZN(g25065) );
NAND2_X4 U_g25066 ( .A1(g23984), .A2(g7195), .ZN(g25066) );
NAND2_X4 U_g25068 ( .A1(g23803), .A2(g5556), .ZN(g25068) );
NAND2_X4 U_g25069 ( .A1(g24014), .A2(g7303), .ZN(g25069) );
NAND2_X4 U_g25070 ( .A1(g24014), .A2(g7391), .ZN(g25070) );
NAND2_X4 U_g25071 ( .A1(g23984), .A2(g7053), .ZN(g25071) );
NAND2_X4 U_g25072 ( .A1(g24014), .A2(g7303), .ZN(g25072) );
NAND2_X4 U_g25073 ( .A1(g24014), .A2(g7391), .ZN(g25073) );
NAND2_X4 U_g25074 ( .A1(g24014), .A2(g7303), .ZN(g25074) );
NAND2_X4 U_g25088 ( .A1(g23950), .A2(g679), .ZN(g25088) );
NAND2_X4 U_g25096 ( .A1(g23979), .A2(g1365), .ZN(g25096) );
NAND2_X4 U_g25106 ( .A1(g24009), .A2(g2059), .ZN(g25106) );
NAND2_X4 U_g25112 ( .A1(g24043), .A2(g2753), .ZN(g25112) );
NAND2_X4 U_g25200 ( .A1(g24965), .A2(g3306), .ZN(g25200) );
NAND2_X4 U_g25203 ( .A1(g24978), .A2(g3462), .ZN(g25203) );
NAND2_X4 U_g25205 ( .A1(g24989), .A2(g3618), .ZN(g25205) );
NAND2_X4 U_g25210 ( .A1(g25000), .A2(g3774), .ZN(g25210) );
NAND4_X4 U_g25312 ( .A1(g21211), .A2(g14442), .A3(g10694), .A4(g24590), .ZN(g25312) );
NAND4_X4 U_g25320 ( .A1(g21219), .A2(g14529), .A3(g10714), .A4(g24595), .ZN(g25320) );
NAND4_X4 U_g25331 ( .A1(g21230), .A2(g14584), .A3(g10735), .A4(g24603), .ZN(g25331) );
NAND4_X4 U_g25340 ( .A1(g21235), .A2(g14618), .A3(g10754), .A4(g24610), .ZN(g25340) );
NAND2_X4 U_g25927 ( .A1(g24965), .A2(g6448), .ZN(g25927) );
NAND2_X4 U_g25928 ( .A1(g24965), .A2(g5438), .ZN(g25928) );
NAND2_X4 U_g25929 ( .A1(g24978), .A2(g6713), .ZN(g25929) );
NAND2_X4 U_g25930 ( .A1(g24978), .A2(g5473), .ZN(g25930) );
NAND2_X4 U_g25931 ( .A1(g24989), .A2(g7015), .ZN(g25931) );
NAND2_X4 U_g25933 ( .A1(g24989), .A2(g5512), .ZN(g25933) );
NAND2_X4 U_g25934 ( .A1(g25000), .A2(g7265), .ZN(g25934) );
NAND2_X4 U_g25936 ( .A1(g25000), .A2(g5556), .ZN(g25936) );
NAND2_X4 U_g25954 ( .A1(g22806), .A2(g24517), .ZN(g25954) );
NAND2_X4 U_g25958 ( .A1(g22847), .A2(g24530), .ZN(g25958) );
NAND2_X4 U_g25964 ( .A1(g22882), .A2(g24543), .ZN(g25964) );
NAND2_X4 U_g25969 ( .A1(g22917), .A2(g24555), .ZN(g25969) );
NAND3_X4 U_g26059 ( .A1(g25422), .A2(g25379), .A3(g25274), .ZN(g26059) );
NAND3_X4 U_g26066 ( .A1(g25431), .A2(g25395), .A3(g25283), .ZN(g26066) );
NAND3_X4 U_g26073 ( .A1(g25438), .A2(g25405), .A3(g25291), .ZN(g26073) );
NAND3_X4 U_g26079 ( .A1(g25445), .A2(g25413), .A3(g25301), .ZN(g26079) );
NAND2_X4 U_g26106 ( .A1(g23644), .A2(g25354), .ZN(g26106) );
NAND4_X4 U_g26119 ( .A1(g8278), .A2(g14657), .A3(g25422), .A4(g25379), .ZN(g26119) );
NAND2_X4 U_g26120 ( .A1(g23694), .A2(g25369), .ZN(g26120) );
NAND4_X4 U_g26129 ( .A1(g8287), .A2(g14691), .A3(g25431), .A4(g25395), .ZN(g26129) );
NAND2_X4 U_g26130 ( .A1(g23748), .A2(g25386), .ZN(g26130) );
NAND4_X4 U_g26143 ( .A1(g8296), .A2(g14725), .A3(g25438), .A4(g25405), .ZN(g26143) );
NAND2_X4 U_g26144 ( .A1(g23803), .A2(g25402), .ZN(g26144) );
NAND4_X4 U_g26148 ( .A1(g8305), .A2(g14753), .A3(g25445), .A4(g25413), .ZN(g26148) );
NAND2_X4 U_g26356 ( .A1(g16539), .A2(g25183), .ZN(g26356) );
NAND2_X4 U_g26399 ( .A1(g16571), .A2(g25186), .ZN(g26399) );
NAND2_X4 U_g26440 ( .A1(g16595), .A2(g25190), .ZN(g26440) );
NAND2_X4 U_g26458 ( .A1(g25343), .A2(g65), .ZN(g26458) );
NAND2_X4 U_g26472 ( .A1(g16615), .A2(g25195), .ZN(g26472) );
NAND2_X4 U_g26482 ( .A1(g25357), .A2(g753), .ZN(g26482) );
NAND2_X4 U_g26498 ( .A1(g25372), .A2(g1439), .ZN(g26498) );
NAND2_X4 U_g26513 ( .A1(g25389), .A2(g2133), .ZN(g26513) );
NAND2_X4 U_g26772 ( .A1(g26320), .A2(g3306), .ZN(g26772) );
NAND2_X4 U_g26779 ( .A1(g26367), .A2(g3462), .ZN(g26779) );
NAND2_X4 U_g26785 ( .A1(g26410), .A2(g3618), .ZN(g26785) );
NAND2_X4 U_g26792 ( .A1(g26451), .A2(g3774), .ZN(g26792) );
NAND2_X4 U_I35020 ( .A1(g26110), .A2(g26099), .ZN(I35020) );
NAND2_X4 U_I35021 ( .A1(g26110), .A2(I35020), .ZN(I35021) );
NAND2_X4 U_I35022 ( .A1(g26099), .A2(I35020), .ZN(I35022) );
NAND2_X4 U_g26859 ( .A1(I35021), .A2(I35022), .ZN(g26859) );
NAND2_X4 U_I35034 ( .A1(g26087), .A2(g26154), .ZN(I35034) );
NAND2_X4 U_I35035 ( .A1(g26087), .A2(I35034), .ZN(I35035) );
NAND2_X4 U_I35036 ( .A1(g26154), .A2(I35034), .ZN(I35036) );
NAND2_X4 U_g26865 ( .A1(I35035), .A2(I35036), .ZN(g26865) );
NAND2_X4 U_I35042 ( .A1(g26151), .A2(g26145), .ZN(I35042) );
NAND2_X4 U_I35043 ( .A1(g26151), .A2(I35042), .ZN(I35043) );
NAND2_X4 U_I35044 ( .A1(g26145), .A2(I35042), .ZN(I35044) );
NAND2_X4 U_g26867 ( .A1(I35043), .A2(I35044), .ZN(g26867) );
NAND2_X4 U_I35057 ( .A1(g26137), .A2(g26126), .ZN(I35057) );
NAND2_X4 U_I35058 ( .A1(g26137), .A2(I35057), .ZN(I35058) );
NAND2_X4 U_I35059 ( .A1(g26126), .A2(I35057), .ZN(I35059) );
NAND2_X4 U_g26874 ( .A1(I35058), .A2(I35059), .ZN(g26874) );
NAND4_X4 U_g26892 ( .A1(g25699), .A2(g26283), .A3(g25569), .A4(g25631), .ZN(g26892) );
NAND3_X4 U_g26902 ( .A1(g25631), .A2(g26283), .A3(g25569), .ZN(g26902) );
NAND4_X4 U_g26906 ( .A1(g25772), .A2(g26327), .A3(g25648), .A4(g25708), .ZN(g26906) );
NAND2_X4 U_g26911 ( .A1(g25569), .A2(g26283), .ZN(g26911) );
NAND3_X4 U_g26915 ( .A1(g25708), .A2(g26327), .A3(g25648), .ZN(g26915) );
NAND4_X4 U_g26918 ( .A1(g25826), .A2(g26374), .A3(g25725), .A4(g25781), .ZN(g26918) );
NAND2_X4 U_g26925 ( .A1(g25648), .A2(g26327), .ZN(g26925) );
NAND3_X4 U_g26928 ( .A1(g25781), .A2(g26374), .A3(g25725), .ZN(g26928) );
NAND4_X4 U_g26931 ( .A1(g25861), .A2(g26417), .A3(g25798), .A4(g25835), .ZN(g26931) );
NAND2_X4 U_I35123 ( .A1(g26107), .A2(g26096), .ZN(I35123) );
NAND2_X4 U_I35124 ( .A1(g26107), .A2(I35123), .ZN(I35124) );
NAND2_X4 U_I35125 ( .A1(g26096), .A2(I35123), .ZN(I35125) );
NAND2_X4 U_g26934 ( .A1(I35124), .A2(I35125), .ZN(g26934) );
NAND2_X4 U_g26938 ( .A1(g25725), .A2(g26374), .ZN(g26938) );
NAND3_X4 U_g26941 ( .A1(g25835), .A2(g26417), .A3(g25798), .ZN(g26941) );
NAND2_X4 U_g26947 ( .A1(g25798), .A2(g26417), .ZN(g26947) );
NAND2_X4 U_g27117 ( .A1(g26320), .A2(g6448), .ZN(g27117) );
NAND2_X4 U_g27118 ( .A1(g26320), .A2(g5438), .ZN(g27118) );
NAND2_X4 U_g27119 ( .A1(g26367), .A2(g6713), .ZN(g27119) );
NAND2_X4 U_g27121 ( .A1(g26367), .A2(g5473), .ZN(g27121) );
NAND2_X4 U_g27122 ( .A1(g26410), .A2(g7015), .ZN(g27122) );
NAND2_X4 U_g27124 ( .A1(g26410), .A2(g5512), .ZN(g27124) );
NAND2_X4 U_g27125 ( .A1(g26451), .A2(g7265), .ZN(g27125) );
NAND2_X4 U_g27130 ( .A1(g26451), .A2(g5556), .ZN(g27130) );
NAND2_X4 U_I35701 ( .A1(g26867), .A2(g26874), .ZN(I35701) );
NAND2_X4 U_I35702 ( .A1(g26867), .A2(I35701), .ZN(I35702) );
NAND2_X4 U_I35703 ( .A1(g26874), .A2(I35701), .ZN(I35703) );
NAND2_X4 U_g27379 ( .A1(I35702), .A2(I35703), .ZN(g27379) );
NAND2_X4 U_I35714 ( .A1(g26859), .A2(g26865), .ZN(I35714) );
NAND2_X4 U_I35715 ( .A1(g26859), .A2(I35714), .ZN(I35715) );
NAND2_X4 U_I35716 ( .A1(g26865), .A2(I35714), .ZN(I35716) );
NAND2_X4 U_g27382 ( .A1(I35715), .A2(I35716), .ZN(g27382) );
NAND2_X4 U_g27390 ( .A1(g26989), .A2(g6448), .ZN(g27390) );
NAND2_X4 U_g27395 ( .A1(g26989), .A2(g5438), .ZN(g27395) );
NAND2_X4 U_g27400 ( .A1(g27012), .A2(g6713), .ZN(g27400) );
NAND2_X4 U_g27408 ( .A1(g27012), .A2(g5473), .ZN(g27408) );
NAND2_X4 U_g27413 ( .A1(g27038), .A2(g7015), .ZN(g27413) );
NAND2_X4 U_g27426 ( .A1(g27038), .A2(g5512), .ZN(g27426) );
NAND2_X4 U_g27431 ( .A1(g27066), .A2(g7265), .ZN(g27431) );
NAND2_X4 U_g27447 ( .A1(g27066), .A2(g5556), .ZN(g27447) );
NAND2_X4 U_I35904 ( .A1(g27051), .A2(g14831), .ZN(I35904) );
NAND2_X4 U_I35905 ( .A1(g27051), .A2(I35904), .ZN(I35905) );
NAND2_X4 U_I35906 ( .A1(g14831), .A2(I35904), .ZN(I35906) );
NAND2_X4 U_g27528 ( .A1(I35905), .A2(I35906), .ZN(g27528) );
NAND2_X4 U_I35944 ( .A1(g27078), .A2(g14904), .ZN(I35944) );
NAND2_X4 U_I35945 ( .A1(g27078), .A2(I35944), .ZN(I35945) );
NAND2_X4 U_I35946 ( .A1(g14904), .A2(I35944), .ZN(I35946) );
NAND2_X4 U_g27550 ( .A1(I35945), .A2(I35946), .ZN(g27550) );
NAND2_X4 U_I35974 ( .A1(g27094), .A2(g14985), .ZN(I35974) );
NAND2_X4 U_I35975 ( .A1(g27094), .A2(I35974), .ZN(I35975) );
NAND2_X4 U_I35976 ( .A1(g14985), .A2(I35974), .ZN(I35976) );
NAND2_X4 U_g27566 ( .A1(I35975), .A2(I35976), .ZN(g27566) );
NAND2_X4 U_g27571 ( .A1(g26869), .A2(g56), .ZN(g27571) );
NAND2_X4 U_I35992 ( .A1(g27106), .A2(g15074), .ZN(I35992) );
NAND2_X4 U_I35993 ( .A1(g27106), .A2(I35992), .ZN(I35993) );
NAND2_X4 U_I35994 ( .A1(g15074), .A2(I35992), .ZN(I35994) );
NAND2_X4 U_g27576 ( .A1(I35993), .A2(I35994), .ZN(g27576) );
NAND2_X4 U_g27580 ( .A1(g26878), .A2(g744), .ZN(g27580) );
NAND2_X4 U_g27583 ( .A1(g26887), .A2(g1430), .ZN(g27583) );
NAND2_X4 U_g27587 ( .A1(g26897), .A2(g2124), .ZN(g27587) );
NAND2_X4 U_g27626 ( .A1(g26989), .A2(g3306), .ZN(g27626) );
NAND2_X4 U_g27627 ( .A1(g27012), .A2(g3462), .ZN(g27627) );
NAND2_X4 U_g27628 ( .A1(g27038), .A2(g3618), .ZN(g27628) );
NAND2_X4 U_g27630 ( .A1(g27066), .A2(g3774), .ZN(g27630) );
NAND2_X4 U_g27738 ( .A1(g25367), .A2(g27415), .ZN(g27738) );
NAND2_X4 U_g27743 ( .A1(g25384), .A2(g27436), .ZN(g27743) );
NAND2_X4 U_g27751 ( .A1(g25400), .A2(g27455), .ZN(g27751) );
NAND2_X4 U_g27756 ( .A1(g25410), .A2(g27471), .ZN(g27756) );
NAND2_X4 U_I36256 ( .A1(g27527), .A2(g15859), .ZN(I36256) );
NAND2_X4 U_I36257 ( .A1(g27527), .A2(I36256), .ZN(I36257) );
NAND2_X4 U_I36258 ( .A1(g15859), .A2(I36256), .ZN(I36258) );
NAND2_X4 U_g27801 ( .A1(I36257), .A2(I36258), .ZN(g27801) );
NAND2_X4 U_I36270 ( .A1(g27549), .A2(g15890), .ZN(I36270) );
NAND2_X4 U_I36271 ( .A1(g27549), .A2(I36270), .ZN(I36271) );
NAND2_X4 U_I36272 ( .A1(g15890), .A2(I36270), .ZN(I36272) );
NAND2_X4 U_g27809 ( .A1(I36271), .A2(I36272), .ZN(g27809) );
NAND2_X4 U_I36289 ( .A1(g27565), .A2(g15923), .ZN(I36289) );
NAND2_X4 U_I36290 ( .A1(g27565), .A2(I36289), .ZN(I36290) );
NAND2_X4 U_I36291 ( .A1(g15923), .A2(I36289), .ZN(I36291) );
NAND2_X4 U_g27830 ( .A1(I36290), .A2(I36291), .ZN(g27830) );
NAND2_X4 U_I36300 ( .A1(g27382), .A2(g27379), .ZN(I36300) );
NAND2_X4 U_I36301 ( .A1(g27382), .A2(I36300), .ZN(I36301) );
NAND2_X4 U_I36302 ( .A1(g27379), .A2(I36300), .ZN(I36302) );
NAND2_X4 U_g27838 ( .A1(I36301), .A2(I36302), .ZN(g27838) );
NAND2_X4 U_I36314 ( .A1(g27575), .A2(g15952), .ZN(I36314) );
NAND2_X4 U_I36315 ( .A1(g27575), .A2(I36314), .ZN(I36315) );
NAND2_X4 U_I36316 ( .A1(g15952), .A2(I36314), .ZN(I36316) );
NAND2_X4 U_g27846 ( .A1(I36315), .A2(I36316), .ZN(g27846) );
NAND2_X4 U_I36591 ( .A1(g27529), .A2(g14885), .ZN(I36591) );
NAND2_X4 U_I36592 ( .A1(g27529), .A2(I36591), .ZN(I36592) );
NAND2_X4 U_I36593 ( .A1(g14885), .A2(I36591), .ZN(I36593) );
NAND2_X4 U_g28046 ( .A1(I36592), .A2(I36593), .ZN(g28046) );
NAND2_X4 U_I36666 ( .A1(g27551), .A2(g14966), .ZN(I36666) );
NAND2_X4 U_I36667 ( .A1(g27551), .A2(I36666), .ZN(I36667) );
NAND2_X4 U_I36668 ( .A1(g14966), .A2(I36666), .ZN(I36668) );
NAND2_X4 U_g28075 ( .A1(I36667), .A2(I36668), .ZN(g28075) );
NAND2_X4 U_I36731 ( .A1(g27567), .A2(g15055), .ZN(I36731) );
NAND2_X4 U_I36732 ( .A1(g27567), .A2(I36731), .ZN(I36732) );
NAND2_X4 U_I36733 ( .A1(g15055), .A2(I36731), .ZN(I36733) );
NAND2_X4 U_g28100 ( .A1(I36732), .A2(I36733), .ZN(g28100) );
NAND2_X4 U_I36779 ( .A1(g27577), .A2(g15151), .ZN(I36779) );
NAND2_X4 U_I36780 ( .A1(g27577), .A2(I36779), .ZN(I36780) );
NAND2_X4 U_I36781 ( .A1(g15151), .A2(I36779), .ZN(I36781) );
NAND2_X4 U_g28118 ( .A1(I36780), .A2(I36781), .ZN(g28118) );
NAND2_X4 U_I37295 ( .A1(g27827), .A2(g27814), .ZN(I37295) );
NAND2_X4 U_I37296 ( .A1(g27827), .A2(I37295), .ZN(I37296) );
NAND2_X4 U_I37297 ( .A1(g27814), .A2(I37295), .ZN(I37297) );
NAND2_X4 U_g28384 ( .A1(I37296), .A2(I37297), .ZN(g28384) );
NAND2_X4 U_I37303 ( .A1(g27802), .A2(g27900), .ZN(I37303) );
NAND2_X4 U_I37304 ( .A1(g27802), .A2(I37303), .ZN(I37304) );
NAND2_X4 U_I37305 ( .A1(g27900), .A2(I37303), .ZN(I37305) );
NAND2_X4 U_g28386 ( .A1(I37304), .A2(I37305), .ZN(g28386) );
NAND2_X4 U_I37311 ( .A1(g27897), .A2(g27883), .ZN(I37311) );
NAND2_X4 U_I37312 ( .A1(g27897), .A2(I37311), .ZN(I37312) );
NAND2_X4 U_I37313 ( .A1(g27883), .A2(I37311), .ZN(I37313) );
NAND2_X4 U_g28388 ( .A1(I37312), .A2(I37313), .ZN(g28388) );
NAND2_X4 U_I37322 ( .A1(g27865), .A2(g27855), .ZN(I37322) );
NAND2_X4 U_I37323 ( .A1(g27865), .A2(I37322), .ZN(I37323) );
NAND2_X4 U_I37324 ( .A1(g27855), .A2(I37322), .ZN(I37324) );
NAND2_X4 U_g28391 ( .A1(I37323), .A2(I37324), .ZN(g28391) );
NAND2_X4 U_I37356 ( .A1(g27824), .A2(g27811), .ZN(I37356) );
NAND2_X4 U_I37357 ( .A1(g27824), .A2(I37356), .ZN(I37357) );
NAND2_X4 U_I37358 ( .A1(g27811), .A2(I37356), .ZN(I37358) );
NAND2_X4 U_g28415 ( .A1(I37357), .A2(I37358), .ZN(g28415) );
NAND2_X4 U_I37813 ( .A1(g28388), .A2(g28391), .ZN(I37813) );
NAND2_X4 U_I37814 ( .A1(g28388), .A2(I37813), .ZN(I37814) );
NAND2_X4 U_I37815 ( .A1(g28391), .A2(I37813), .ZN(I37815) );
NAND2_X4 U_g28842 ( .A1(I37814), .A2(I37815), .ZN(g28842) );
NAND2_X4 U_I37822 ( .A1(g28384), .A2(g28386), .ZN(I37822) );
NAND2_X4 U_I37823 ( .A1(g28384), .A2(I37822), .ZN(I37823) );
NAND2_X4 U_I37824 ( .A1(g28386), .A2(I37822), .ZN(I37824) );
NAND2_X4 U_g28845 ( .A1(I37823), .A2(I37824), .ZN(g28845) );
NAND2_X4 U_g28978 ( .A1(g9150), .A2(g28512), .ZN(g28978) );
NAND2_X4 U_g29001 ( .A1(g9161), .A2(g28512), .ZN(g29001) );
NAND2_X4 U_g29008 ( .A1(g9174), .A2(g28540), .ZN(g29008) );
NAND2_X4 U_g29026 ( .A1(g9187), .A2(g28512), .ZN(g29026) );
NAND2_X4 U_g29030 ( .A1(g9203), .A2(g28540), .ZN(g29030) );
NAND2_X4 U_g29038 ( .A1(g9216), .A2(g28567), .ZN(g29038) );
NAND2_X4 U_g29045 ( .A1(g9232), .A2(g28512), .ZN(g29045) );
NAND2_X4 U_g29049 ( .A1(g9248), .A2(g28540), .ZN(g29049) );
NAND2_X4 U_g29053 ( .A1(g9264), .A2(g28567), .ZN(g29053) );
NAND2_X4 U_g29060 ( .A1(g9277), .A2(g28595), .ZN(g29060) );
NAND2_X4 U_g29062 ( .A1(g9310), .A2(g28540), .ZN(g29062) );
NAND2_X4 U_g29068 ( .A1(g9326), .A2(g28567), .ZN(g29068) );
NAND2_X4 U_g29072 ( .A1(g9342), .A2(g28595), .ZN(g29072) );
NAND2_X4 U_g29076 ( .A1(g9391), .A2(g28567), .ZN(g29076) );
NAND2_X4 U_g29080 ( .A1(g9407), .A2(g28595), .ZN(g29080) );
NAND2_X4 U_g29087 ( .A1(g9488), .A2(g28595), .ZN(g29087) );
NAND2_X4 U_g29088 ( .A1(g9507), .A2(g28512), .ZN(g29088) );
NAND2_X4 U_g29096 ( .A1(g9649), .A2(g28540), .ZN(g29096) );
NAND2_X4 U_g29103 ( .A1(g9795), .A2(g28567), .ZN(g29103) );
NAND2_X4 U_g29107 ( .A1(g9941), .A2(g28595), .ZN(g29107) );
NAND2_X4 U_I38378 ( .A1(g28845), .A2(g28842), .ZN(I38378) );
NAND2_X4 U_I38379 ( .A1(g28845), .A2(I38378), .ZN(I38379) );
NAND2_X4 U_I38380 ( .A1(g28842), .A2(I38378), .ZN(I38380) );
NAND2_X4 U_g29265 ( .A1(I38379), .A2(I38380), .ZN(g29265) );
NAND2_X4 U_I38810 ( .A1(g29303), .A2(g15904), .ZN(I38810) );
NAND2_X4 U_I38811 ( .A1(g29303), .A2(I38810), .ZN(I38811) );
NAND2_X4 U_I38812 ( .A1(g15904), .A2(I38810), .ZN(I38812) );
NAND2_X4 U_g29498 ( .A1(I38811), .A2(I38812), .ZN(g29498) );
NAND2_X4 U_I38820 ( .A1(g29313), .A2(g15933), .ZN(I38820) );
NAND2_X4 U_I38821 ( .A1(g29313), .A2(I38820), .ZN(I38821) );
NAND2_X4 U_I38822 ( .A1(g15933), .A2(I38820), .ZN(I38822) );
NAND2_X4 U_g29500 ( .A1(I38821), .A2(I38822), .ZN(g29500) );
NAND2_X4 U_I38831 ( .A1(g29324), .A2(g15962), .ZN(I38831) );
NAND2_X4 U_I38832 ( .A1(g29324), .A2(I38831), .ZN(I38832) );
NAND2_X4 U_I38833 ( .A1(g15962), .A2(I38831), .ZN(I38833) );
NAND2_X4 U_g29503 ( .A1(I38832), .A2(I38833), .ZN(g29503) );
NAND2_X4 U_I38841 ( .A1(g29333), .A2(g15981), .ZN(I38841) );
NAND2_X4 U_I38842 ( .A1(g29333), .A2(I38841), .ZN(I38842) );
NAND2_X4 U_I38843 ( .A1(g15981), .A2(I38841), .ZN(I38843) );
NAND2_X4 U_g29505 ( .A1(I38842), .A2(I38843), .ZN(g29505) );
NAND2_X4 U_I39323 ( .A1(g29721), .A2(g29713), .ZN(I39323) );
NAND2_X4 U_I39324 ( .A1(g29721), .A2(I39323), .ZN(I39324) );
NAND2_X4 U_I39325 ( .A1(g29713), .A2(I39323), .ZN(I39325) );
NAND2_X4 U_g29911 ( .A1(I39324), .A2(I39325), .ZN(g29911) );
NAND2_X4 U_I39331 ( .A1(g29705), .A2(g29751), .ZN(I39331) );
NAND2_X4 U_I39332 ( .A1(g29705), .A2(I39331), .ZN(I39332) );
NAND2_X4 U_I39333 ( .A1(g29751), .A2(I39331), .ZN(I39333) );
NAND2_X4 U_g29913 ( .A1(I39332), .A2(I39333), .ZN(g29913) );
NAND2_X4 U_I39339 ( .A1(g29748), .A2(g29741), .ZN(I39339) );
NAND2_X4 U_I39340 ( .A1(g29748), .A2(I39339), .ZN(I39340) );
NAND2_X4 U_I39341 ( .A1(g29741), .A2(I39339), .ZN(I39341) );
NAND2_X4 U_g29915 ( .A1(I39340), .A2(I39341), .ZN(g29915) );
NAND2_X4 U_I39347 ( .A1(g29732), .A2(g29728), .ZN(I39347) );
NAND2_X4 U_I39348 ( .A1(g29732), .A2(I39347), .ZN(I39348) );
NAND2_X4 U_I39349 ( .A1(g29728), .A2(I39347), .ZN(I39349) );
NAND2_X4 U_g29917 ( .A1(I39348), .A2(I39349), .ZN(g29917) );
NAND2_X4 U_I39359 ( .A1(g29766), .A2(g15880), .ZN(I39359) );
NAND2_X4 U_I39360 ( .A1(g29766), .A2(I39359), .ZN(I39360) );
NAND2_X4 U_I39361 ( .A1(g15880), .A2(I39359), .ZN(I39361) );
NAND2_X4 U_g29923 ( .A1(I39360), .A2(I39361), .ZN(g29923) );
NAND2_X4 U_I39367 ( .A1(g29767), .A2(g15913), .ZN(I39367) );
NAND2_X4 U_I39368 ( .A1(g29767), .A2(I39367), .ZN(I39368) );
NAND2_X4 U_I39369 ( .A1(g15913), .A2(I39367), .ZN(I39369) );
NAND2_X4 U_g29925 ( .A1(I39368), .A2(I39369), .ZN(g29925) );
NAND2_X4 U_I39375 ( .A1(g29768), .A2(g15942), .ZN(I39375) );
NAND2_X4 U_I39376 ( .A1(g29768), .A2(I39375), .ZN(I39376) );
NAND2_X4 U_I39377 ( .A1(g15942), .A2(I39375), .ZN(I39377) );
NAND2_X4 U_g29927 ( .A1(I39376), .A2(I39377), .ZN(g29927) );
NAND2_X4 U_I39384 ( .A1(g29718), .A2(g29710), .ZN(I39384) );
NAND2_X4 U_I39385 ( .A1(g29718), .A2(I39384), .ZN(I39385) );
NAND2_X4 U_I39386 ( .A1(g29710), .A2(I39384), .ZN(I39386) );
NAND2_X4 U_g29930 ( .A1(I39385), .A2(I39386), .ZN(g29930) );
NAND2_X4 U_I39391 ( .A1(g29769), .A2(g15971), .ZN(I39391) );
NAND2_X4 U_I39392 ( .A1(g29769), .A2(I39391), .ZN(I39392) );
NAND2_X4 U_I39393 ( .A1(g15971), .A2(I39391), .ZN(I39393) );
NAND2_X4 U_g29931 ( .A1(I39392), .A2(I39393), .ZN(g29931) );
NAND2_X4 U_I39532 ( .A1(g29915), .A2(g29917), .ZN(I39532) );
NAND2_X4 U_I39533 ( .A1(g29915), .A2(I39532), .ZN(I39533) );
NAND2_X4 U_I39534 ( .A1(g29917), .A2(I39532), .ZN(I39534) );
NAND2_X4 U_g30034 ( .A1(I39533), .A2(I39534), .ZN(g30034) );
NAND2_X4 U_I39539 ( .A1(g29911), .A2(g29913), .ZN(I39539) );
NAND2_X4 U_I39540 ( .A1(g29911), .A2(I39539), .ZN(I39540) );
NAND2_X4 U_I39541 ( .A1(g29913), .A2(I39539), .ZN(I39541) );
NAND2_X4 U_g30035 ( .A1(I39540), .A2(I39541), .ZN(g30035) );
NAND2_X4 U_I39689 ( .A1(g30035), .A2(g30034), .ZN(I39689) );
NAND2_X4 U_I39690 ( .A1(g30035), .A2(I39689), .ZN(I39690) );
NAND2_X4 U_I39691 ( .A1(g30034), .A2(I39689), .ZN(I39691) );
NAND2_X4 U_g30228 ( .A1(I39690), .A2(I39691), .ZN(g30228) );
NAND2_X4 U_I40558 ( .A1(g30605), .A2(g30597), .ZN(I40558) );
NAND2_X4 U_I40559 ( .A1(g30605), .A2(I40558), .ZN(I40559) );
NAND2_X4 U_I40560 ( .A1(g30597), .A2(I40558), .ZN(I40560) );
NAND2_X4 U_g30768 ( .A1(I40559), .A2(I40560), .ZN(g30768) );
NAND2_X4 U_I40571 ( .A1(g30588), .A2(g30632), .ZN(I40571) );
NAND2_X4 U_I40572 ( .A1(g30588), .A2(I40571), .ZN(I40572) );
NAND2_X4 U_I40573 ( .A1(g30632), .A2(I40571), .ZN(I40573) );
NAND2_X4 U_g30771 ( .A1(I40572), .A2(I40573), .ZN(g30771) );
NAND2_X4 U_I40587 ( .A1(g30629), .A2(g30622), .ZN(I40587) );
NAND2_X4 U_I40588 ( .A1(g30629), .A2(I40587), .ZN(I40588) );
NAND2_X4 U_I40589 ( .A1(g30622), .A2(I40587), .ZN(I40589) );
NAND2_X4 U_g30775 ( .A1(I40588), .A2(I40589), .ZN(g30775) );
NAND2_X4 U_I40603 ( .A1(g30614), .A2(g30610), .ZN(I40603) );
NAND2_X4 U_I40604 ( .A1(g30614), .A2(I40603), .ZN(I40604) );
NAND2_X4 U_I40605 ( .A1(g30610), .A2(I40603), .ZN(I40605) );
NAND2_X4 U_g30779 ( .A1(I40604), .A2(I40605), .ZN(g30779) );
NAND2_X4 U_I40627 ( .A1(g30602), .A2(g30594), .ZN(I40627) );
NAND2_X4 U_I40628 ( .A1(g30602), .A2(I40627), .ZN(I40628) );
NAND2_X4 U_I40629 ( .A1(g30594), .A2(I40627), .ZN(I40629) );
NAND2_X4 U_g30791 ( .A1(I40628), .A2(I40629), .ZN(g30791) );
NAND2_X4 U_I41010 ( .A1(g30775), .A2(g30779), .ZN(I41010) );
NAND2_X4 U_I41011 ( .A1(g30775), .A2(I41010), .ZN(I41011) );
NAND2_X4 U_I41012 ( .A1(g30779), .A2(I41010), .ZN(I41012) );
NAND2_X4 U_g30926 ( .A1(I41011), .A2(I41012), .ZN(g30926) );
NAND2_X4 U_I41017 ( .A1(g30768), .A2(g30771), .ZN(I41017) );
NAND2_X4 U_I41018 ( .A1(g30768), .A2(I41017), .ZN(I41018) );
NAND2_X4 U_I41019 ( .A1(g30771), .A2(I41017), .ZN(I41019) );
NAND2_X4 U_g30927 ( .A1(I41018), .A2(I41019), .ZN(g30927) );
NAND2_X4 U_I41064 ( .A1(g30927), .A2(g30926), .ZN(I41064) );
NAND2_X4 U_I41065 ( .A1(g30927), .A2(I41064), .ZN(I41065) );
NAND2_X4 U_I41066 ( .A1(g30926), .A2(I41064), .ZN(I41066) );
NAND2_X4 U_g30952 ( .A1(I41065), .A2(I41066), .ZN(g30952) );
NOR3_X4 U_g7528 ( .A1(g3151), .A2(g3142), .A3(g3147), .ZN(g7528) );
NOR2_X4 U_g7575 ( .A1(g2984), .A2(g2985), .ZN(g7575) );
NOR2_X4 U_g7795 ( .A1(g2992), .A2(g2991), .ZN(g7795) );
NOR4_X4 U_g8430 ( .A1(g3198), .A2(g8120), .A3(g3194), .A4(g3191), .ZN(g8430) );
NOR3_X4 U_g10784 ( .A1(g5630), .A2(g5649), .A3(g5676), .ZN(g10784) );
NOR3_X4 U_g10789 ( .A1(g5650), .A2(g5677), .A3(g5709), .ZN(g10789) );
NOR3_X4 U_g10793 ( .A1(g5658), .A2(g5687), .A3(g5728), .ZN(g10793) );
NOR3_X4 U_g10797 ( .A1(g5678), .A2(g5710), .A3(g5757), .ZN(g10797) );
NOR3_X4 U_g10801 ( .A1(g5688), .A2(g5729), .A3(g5767), .ZN(g10801) );
NOR3_X4 U_g10805 ( .A1(g5696), .A2(g5739), .A3(g5786), .ZN(g10805) );
NOR3_X4 U_g10810 ( .A1(g5711), .A2(g5758), .A3(g5807), .ZN(g10810) );
NOR3_X4 U_g10814 ( .A1(g5730), .A2(g5768), .A3(g5816), .ZN(g10814) );
NOR3_X4 U_g10818 ( .A1(g5740), .A2(g5787), .A3(g5826), .ZN(g10818) );
NOR3_X4 U_g10822 ( .A1(g5748), .A2(g5797), .A3(g5845), .ZN(g10822) );
NOR3_X4 U_g10831 ( .A1(g5769), .A2(g5817), .A3(g5863), .ZN(g10831) );
NOR3_X4 U_g10835 ( .A1(g5788), .A2(g5827), .A3(g5872), .ZN(g10835) );
NOR3_X4 U_g10839 ( .A1(g5798), .A2(g5846), .A3(g5882), .ZN(g10839) );
NOR3_X4 U_g10851 ( .A1(g5828), .A2(g5873), .A3(g5910), .ZN(g10851) );
NOR3_X4 U_g10855 ( .A1(g5847), .A2(g5883), .A3(g5919), .ZN(g10855) );
NOR3_X4 U_g10872 ( .A1(g5884), .A2(g5920), .A3(g5949), .ZN(g10872) );
NOR3_X4 U_g11600 ( .A1(g9049), .A2(g9064), .A3(g9078), .ZN(g11600) );
NOR4_X4 U_g11622 ( .A1(g8183), .A2(g11332), .A3(g7928), .A4(g11069), .ZN(g11622) );
NOR3_X4 U_g11624 ( .A1(g9062), .A2(g9075), .A3(g9091), .ZN(g11624) );
NOR3_X4 U_g11627 ( .A1(g9063), .A2(g9077), .A3(g9093), .ZN(g11627) );
NOR3_X4 U_g11630 ( .A1(g9066), .A2(g9081), .A3(g9097), .ZN(g11630) );
NOR4_X4 U_g11643 ( .A1(g11481), .A2(g8045), .A3(g7928), .A4(g11069), .ZN(g11643) );
NOR3_X4 U_g11644 ( .A1(g9076), .A2(g9092), .A3(g9102), .ZN(g11644) );
NOR3_X4 U_g11647 ( .A1(g9079), .A2(g9094), .A3(g9103), .ZN(g11647) );
NOR3_X4 U_g11650 ( .A1(g9080), .A2(g9096), .A3(g9105), .ZN(g11650) );
NOR3_X4 U_g11653 ( .A1(g9083), .A2(g9100), .A3(g9109), .ZN(g11653) );
NOR4_X4 U_g11660 ( .A1(g8183), .A2(g8045), .A3(g7928), .A4(g11069), .ZN(g11660) );
NOR3_X4 U_g11663 ( .A1(g9095), .A2(g9104), .A3(g9112), .ZN(g11663) );
NOR3_X4 U_g11666 ( .A1(g9098), .A2(g9106), .A3(g9113), .ZN(g11666) );
NOR3_X4 U_g11669 ( .A1(g9099), .A2(g9108), .A3(g9115), .ZN(g11669) );
NOR3_X4 U_g11675 ( .A1(g9107), .A2(g9114), .A3(g9120), .ZN(g11675) );
NOR3_X4 U_g11678 ( .A1(g9110), .A2(g9116), .A3(g9121), .ZN(g11678) );
NOR3_X4 U_g11681 ( .A1(g9111), .A2(g9118), .A3(g9123), .ZN(g11681) );
NOR3_X4 U_g11687 ( .A1(g9117), .A2(g9122), .A3(g9126), .ZN(g11687) );
NOR3_X4 U_g11690 ( .A1(g9119), .A2(g9124), .A3(g9127), .ZN(g11690) );
NOR3_X4 U_g11697 ( .A1(g9125), .A2(g9131), .A3(g9133), .ZN(g11697) );
NOR3_X4 U_g11703 ( .A1(g9132), .A2(g9137), .A3(g9139), .ZN(g11703) );
NOR3_X4 U_g11711 ( .A1(g9138), .A2(g9143), .A3(g9145), .ZN(g11711) );
NOR3_X4 U_g11744 ( .A1(g9241), .A2(g9301), .A3(g9364), .ZN(g11744) );
NOR3_X4 U_g11759 ( .A1(g9302), .A2(g9365), .A3(g9438), .ZN(g11759) );
NOR3_X4 U_g11760 ( .A1(g9319), .A2(g9382), .A3(g9461), .ZN(g11760) );
NOR3_X4 U_g11767 ( .A1(g9366), .A2(g9439), .A3(g9518), .ZN(g11767) );
NOR3_X4 U_g11768 ( .A1(g9367), .A2(g9441), .A3(g9521), .ZN(g11768) );
NOR3_X4 U_g11772 ( .A1(g9383), .A2(g9462), .A3(g9580), .ZN(g11772) );
NOR3_X4 U_g11773 ( .A1(g9400), .A2(g9479), .A3(g9603), .ZN(g11773) );
NOR3_X4 U_g11780 ( .A1(g9440), .A2(g9519), .A3(g9630), .ZN(g11780) );
NOR3_X4 U_g11781 ( .A1(g9442), .A2(g9522), .A3(g9633), .ZN(g11781) );
NOR3_X4 U_g11784 ( .A1(g9463), .A2(g9581), .A3(g9660), .ZN(g11784) );
NOR3_X4 U_g11785 ( .A1(g9464), .A2(g9583), .A3(g9663), .ZN(g11785) );
NOR3_X4 U_g11789 ( .A1(g9480), .A2(g9604), .A3(g9722), .ZN(g11789) );
NOR3_X4 U_g11790 ( .A1(g9497), .A2(g9621), .A3(g9745), .ZN(g11790) );
NOR3_X4 U_g11799 ( .A1(g9520), .A2(g9631), .A3(g9759), .ZN(g11799) );
NOR3_X4 U_g11800 ( .A1(g9523), .A2(g9634), .A3(g9762), .ZN(g11800) );
NOR3_X4 U_g11806 ( .A1(g9582), .A2(g9661), .A3(g9776), .ZN(g11806) );
NOR3_X4 U_g11807 ( .A1(g9584), .A2(g9664), .A3(g9779), .ZN(g11807) );
NOR3_X4 U_g11810 ( .A1(g9605), .A2(g9723), .A3(g9806), .ZN(g11810) );
NOR3_X4 U_g11811 ( .A1(g9606), .A2(g9725), .A3(g9809), .ZN(g11811) );
NOR3_X4 U_g11815 ( .A1(g9622), .A2(g9746), .A3(g9868), .ZN(g11815) );
NOR3_X4 U_g11822 ( .A1(g9632), .A2(g9760), .A3(g9888), .ZN(g11822) );
NOR3_X4 U_g11823 ( .A1(g9635), .A2(g9763), .A3(g9891), .ZN(g11823) );
NOR3_X4 U_g11828 ( .A1(g9639), .A2(g9764), .A3(g9892), .ZN(g11828) );
NOR3_X4 U_g11830 ( .A1(g9647), .A2(g9773), .A3(g9901), .ZN(g11830) );
NOR3_X4 U_g11831 ( .A1(g9648), .A2(g9775), .A3(g9904), .ZN(g11831) );
NOR3_X4 U_g11832 ( .A1(g9662), .A2(g9777), .A3(g9905), .ZN(g11832) );
NOR3_X4 U_g11833 ( .A1(g9665), .A2(g9780), .A3(g9908), .ZN(g11833) );
NOR3_X4 U_g11839 ( .A1(g9724), .A2(g9807), .A3(g9922), .ZN(g11839) );
NOR3_X4 U_g11840 ( .A1(g9726), .A2(g9810), .A3(g9925), .ZN(g11840) );
NOR3_X4 U_g11843 ( .A1(g9747), .A2(g9869), .A3(g9952), .ZN(g11843) );
NOR3_X4 U_g11844 ( .A1(g9748), .A2(g9871), .A3(g9955), .ZN(g11844) );
NOR3_X4 U_g11855 ( .A1(g9761), .A2(g9889), .A3(g10009), .ZN(g11855) );
NOR3_X4 U_g11860 ( .A1(g9765), .A2(g9893), .A3(g10012), .ZN(g11860) );
NOR3_X4 U_g11861 ( .A1(g9766), .A2(g9894), .A3(g10013), .ZN(g11861) );
NOR3_X4 U_g11863 ( .A1(g9774), .A2(g9902), .A3(g10035), .ZN(g11863) );
NOR3_X4 U_g11864 ( .A1(g9778), .A2(g9906), .A3(g10042), .ZN(g11864) );
NOR3_X4 U_g11865 ( .A1(g9781), .A2(g9909), .A3(g10045), .ZN(g11865) );
NOR3_X4 U_g11870 ( .A1(g9785), .A2(g9910), .A3(g10046), .ZN(g11870) );
NOR3_X4 U_g11872 ( .A1(g9793), .A2(g9919), .A3(g10055), .ZN(g11872) );
NOR3_X4 U_g11873 ( .A1(g9794), .A2(g9921), .A3(g10058), .ZN(g11873) );
NOR3_X4 U_g11874 ( .A1(g9808), .A2(g9923), .A3(g10059), .ZN(g11874) );
NOR3_X4 U_g11875 ( .A1(g9811), .A2(g9926), .A3(g10062), .ZN(g11875) );
NOR3_X4 U_g11881 ( .A1(g9870), .A2(g9953), .A3(g10076), .ZN(g11881) );
NOR3_X4 U_g11882 ( .A1(g9872), .A2(g9956), .A3(g10079), .ZN(g11882) );
NOR3_X4 U_g11889 ( .A1(g9887), .A2(g10007), .A3(g10101), .ZN(g11889) );
NOR3_X4 U_g11890 ( .A1(g9890), .A2(g10010), .A3(g10103), .ZN(g11890) );
NOR3_X4 U_g11896 ( .A1(g9903), .A2(g10036), .A3(g10112), .ZN(g11896) );
NOR3_X4 U_g11897 ( .A1(g9907), .A2(g10043), .A3(g10118), .ZN(g11897) );
NOR3_X4 U_g11902 ( .A1(g9911), .A2(g10047), .A3(g10121), .ZN(g11902) );
NOR3_X4 U_g11903 ( .A1(g9912), .A2(g10048), .A3(g10122), .ZN(g11903) );
NOR3_X4 U_g11905 ( .A1(g9920), .A2(g10056), .A3(g10144), .ZN(g11905) );
NOR3_X4 U_g11906 ( .A1(g9924), .A2(g10060), .A3(g10151), .ZN(g11906) );
NOR3_X4 U_g11907 ( .A1(g9927), .A2(g10063), .A3(g10154), .ZN(g11907) );
NOR3_X4 U_g11912 ( .A1(g9931), .A2(g10064), .A3(g10155), .ZN(g11912) );
NOR3_X4 U_g11914 ( .A1(g9939), .A2(g10073), .A3(g10164), .ZN(g11914) );
NOR3_X4 U_g11915 ( .A1(g9940), .A2(g10075), .A3(g10167), .ZN(g11915) );
NOR3_X4 U_g11916 ( .A1(g9954), .A2(g10077), .A3(g10168), .ZN(g11916) );
NOR3_X4 U_g11917 ( .A1(g9957), .A2(g10080), .A3(g10171), .ZN(g11917) );
NOR3_X4 U_g11928 ( .A1(g10008), .A2(g10102), .A3(g10192), .ZN(g11928) );
NOR3_X4 U_g11934 ( .A1(g10011), .A2(g10104), .A3(g10193), .ZN(g11934) );
NOR3_X4 U_g11935 ( .A1(g10014), .A2(g10106), .A3(g10196), .ZN(g11935) );
NOR3_X4 U_g11938 ( .A1(g10037), .A2(g10113), .A3(g10201), .ZN(g11938) );
NOR3_X4 U_g11939 ( .A1(g10041), .A2(g10116), .A3(g10206), .ZN(g11939) );
NOR3_X4 U_g11940 ( .A1(g10044), .A2(g10119), .A3(g10208), .ZN(g11940) );
NOR3_X4 U_g11946 ( .A1(g10057), .A2(g10145), .A3(g10217), .ZN(g11946) );
NOR3_X4 U_g11947 ( .A1(g10061), .A2(g10152), .A3(g10223), .ZN(g11947) );
NOR3_X4 U_g11952 ( .A1(g10065), .A2(g10156), .A3(g10226), .ZN(g11952) );
NOR3_X4 U_g11953 ( .A1(g10066), .A2(g10157), .A3(g10227), .ZN(g11953) );
NOR3_X4 U_g11955 ( .A1(g10074), .A2(g10165), .A3(g10249), .ZN(g11955) );
NOR3_X4 U_g11956 ( .A1(g10078), .A2(g10169), .A3(g10256), .ZN(g11956) );
NOR3_X4 U_g11957 ( .A1(g10081), .A2(g10172), .A3(g10259), .ZN(g11957) );
NOR3_X4 U_g11962 ( .A1(g10085), .A2(g10173), .A3(g10260), .ZN(g11962) );
NOR3_X4 U_g11964 ( .A1(g10093), .A2(g10182), .A3(g10269), .ZN(g11964) );
NOR3_X4 U_g11965 ( .A1(g10094), .A2(g10184), .A3(g10272), .ZN(g11965) );
NOR3_X4 U_g11974 ( .A1(g10105), .A2(g10194), .A3(g10279), .ZN(g11974) );
NOR3_X4 U_g11975 ( .A1(g10107), .A2(g10197), .A3(g10282), .ZN(g11975) );
NOR3_X4 U_g11979 ( .A1(g10114), .A2(g10202), .A3(g10288), .ZN(g11979) );
NOR3_X4 U_g11980 ( .A1(g10115), .A2(g10204), .A3(g10291), .ZN(g11980) );
NOR3_X4 U_g11981 ( .A1(g10117), .A2(g10207), .A3(g10294), .ZN(g11981) );
NOR3_X4 U_g11987 ( .A1(g10120), .A2(g10209), .A3(g10295), .ZN(g11987) );
NOR3_X4 U_g11988 ( .A1(g10123), .A2(g10211), .A3(g10298), .ZN(g11988) );
NOR3_X4 U_g11991 ( .A1(g10146), .A2(g10218), .A3(g10303), .ZN(g11991) );
NOR3_X4 U_g11992 ( .A1(g10150), .A2(g10221), .A3(g10308), .ZN(g11992) );
NOR3_X4 U_g11993 ( .A1(g10153), .A2(g10224), .A3(g10310), .ZN(g11993) );
NOR3_X4 U_g11999 ( .A1(g10166), .A2(g10250), .A3(g10319), .ZN(g11999) );
NOR3_X4 U_g12000 ( .A1(g10170), .A2(g10257), .A3(g10325), .ZN(g12000) );
NOR3_X4 U_g12005 ( .A1(g10174), .A2(g10261), .A3(g10328), .ZN(g12005) );
NOR3_X4 U_g12006 ( .A1(g10175), .A2(g10262), .A3(g10329), .ZN(g12006) );
NOR3_X4 U_g12008 ( .A1(g10183), .A2(g10270), .A3(g10351), .ZN(g12008) );
NOR3_X4 U_g12026 ( .A1(g10195), .A2(g10280), .A3(g10360), .ZN(g12026) );
NOR3_X4 U_g12033 ( .A1(g10199), .A2(g10284), .A3(g10362), .ZN(g12033) );
NOR3_X4 U_g12034 ( .A1(g10200), .A2(g10286), .A3(g10365), .ZN(g12034) );
NOR3_X4 U_g12035 ( .A1(g10203), .A2(g10289), .A3(g10367), .ZN(g12035) );
NOR3_X4 U_g12036 ( .A1(g10205), .A2(g10292), .A3(g10370), .ZN(g12036) );
NOR3_X4 U_g12043 ( .A1(g10210), .A2(g10296), .A3(g10372), .ZN(g12043) );
NOR3_X4 U_g12044 ( .A1(g10212), .A2(g10299), .A3(g10375), .ZN(g12044) );
NOR3_X4 U_g12048 ( .A1(g10219), .A2(g10304), .A3(g10381), .ZN(g12048) );
NOR3_X4 U_g12049 ( .A1(g10220), .A2(g10306), .A3(g10384), .ZN(g12049) );
NOR3_X4 U_g12050 ( .A1(g10222), .A2(g10309), .A3(g10387), .ZN(g12050) );
NOR3_X4 U_g12056 ( .A1(g10225), .A2(g10311), .A3(g10388), .ZN(g12056) );
NOR3_X4 U_g12057 ( .A1(g10228), .A2(g10313), .A3(g10391), .ZN(g12057) );
NOR3_X4 U_g12060 ( .A1(g10251), .A2(g10320), .A3(g10396), .ZN(g12060) );
NOR3_X4 U_g12061 ( .A1(g10255), .A2(g10323), .A3(g10401), .ZN(g12061) );
NOR3_X4 U_g12062 ( .A1(g10258), .A2(g10326), .A3(g10403), .ZN(g12062) );
NOR3_X4 U_g12068 ( .A1(g10271), .A2(g10352), .A3(g10412), .ZN(g12068) );
NOR3_X4 U_g12079 ( .A1(g10281), .A2(g10361), .A3(g10422), .ZN(g12079) );
NOR3_X4 U_g12080 ( .A1(g10285), .A2(g10363), .A3(g10430), .ZN(g12080) );
NOR3_X4 U_g12081 ( .A1(g10287), .A2(g10366), .A3(g10433), .ZN(g12081) );
NOR3_X4 U_g12082 ( .A1(g10290), .A2(g10368), .A3(g10435), .ZN(g12082) );
NOR3_X4 U_g12083 ( .A1(g10293), .A2(g10371), .A3(g10438), .ZN(g12083) );
NOR3_X4 U_g12090 ( .A1(g10297), .A2(g10373), .A3(g10439), .ZN(g12090) );
NOR3_X4 U_g12097 ( .A1(g10301), .A2(g10377), .A3(g10441), .ZN(g12097) );
NOR3_X4 U_g12098 ( .A1(g10302), .A2(g10379), .A3(g10444), .ZN(g12098) );
NOR3_X4 U_g12099 ( .A1(g10305), .A2(g10382), .A3(g10446), .ZN(g12099) );
NOR3_X4 U_g12100 ( .A1(g10307), .A2(g10385), .A3(g10449), .ZN(g12100) );
NOR3_X4 U_g12107 ( .A1(g10312), .A2(g10389), .A3(g10451), .ZN(g12107) );
NOR3_X4 U_g12108 ( .A1(g10314), .A2(g10392), .A3(g10454), .ZN(g12108) );
NOR3_X4 U_g12112 ( .A1(g10321), .A2(g10397), .A3(g10460), .ZN(g12112) );
NOR3_X4 U_g12113 ( .A1(g10322), .A2(g10399), .A3(g10463), .ZN(g12113) );
NOR3_X4 U_g12114 ( .A1(g10324), .A2(g10402), .A3(g10466), .ZN(g12114) );
NOR3_X4 U_g12120 ( .A1(g10327), .A2(g10404), .A3(g10467), .ZN(g12120) );
NOR3_X4 U_g12121 ( .A1(g10330), .A2(g10406), .A3(g10470), .ZN(g12121) );
NOR3_X4 U_g12124 ( .A1(g10353), .A2(g10413), .A3(g10475), .ZN(g12124) );
NOR3_X4 U_g12145 ( .A1(g10364), .A2(g10431), .A3(g10492), .ZN(g12145) );
NOR3_X4 U_g12146 ( .A1(g10369), .A2(g10436), .A3(g10496), .ZN(g12146) );
NOR3_X4 U_g12151 ( .A1(g10374), .A2(g10440), .A3(g10498), .ZN(g12151) );
NOR3_X4 U_g12152 ( .A1(g10378), .A2(g10442), .A3(g10506), .ZN(g12152) );
NOR3_X4 U_g12153 ( .A1(g10380), .A2(g10445), .A3(g10509), .ZN(g12153) );
NOR3_X4 U_g12154 ( .A1(g10383), .A2(g10447), .A3(g10511), .ZN(g12154) );
NOR3_X4 U_g12155 ( .A1(g10386), .A2(g10450), .A3(g10514), .ZN(g12155) );
NOR3_X4 U_g12162 ( .A1(g10390), .A2(g10452), .A3(g10515), .ZN(g12162) );
NOR3_X4 U_g12169 ( .A1(g10394), .A2(g10456), .A3(g10517), .ZN(g12169) );
NOR3_X4 U_g12170 ( .A1(g10395), .A2(g10458), .A3(g10520), .ZN(g12170) );
NOR3_X4 U_g12171 ( .A1(g10398), .A2(g10461), .A3(g10522), .ZN(g12171) );
NOR3_X4 U_g12172 ( .A1(g10400), .A2(g10464), .A3(g10525), .ZN(g12172) );
NOR3_X4 U_g12179 ( .A1(g10405), .A2(g10468), .A3(g10527), .ZN(g12179) );
NOR3_X4 U_g12180 ( .A1(g10407), .A2(g10471), .A3(g10530), .ZN(g12180) );
NOR3_X4 U_g12184 ( .A1(g10414), .A2(g10476), .A3(g10536), .ZN(g12184) );
NOR3_X4 U_g12185 ( .A1(g10415), .A2(g10478), .A3(g10539), .ZN(g12185) );
NOR3_X4 U_g12192 ( .A1(g10423), .A2(g10485), .A3(g10548), .ZN(g12192) );
NOR3_X4 U_g12193 ( .A1(g10432), .A2(g10493), .A3(g10555), .ZN(g12193) );
NOR3_X4 U_g12194 ( .A1(g10434), .A2(g10494), .A3(g10556), .ZN(g12194) );
NOR3_X4 U_g12195 ( .A1(g10437), .A2(g10497), .A3(g10558), .ZN(g12195) );
NOR3_X4 U_g12207 ( .A1(g10443), .A2(g10507), .A3(g10566), .ZN(g12207) );
NOR3_X4 U_g12208 ( .A1(g10448), .A2(g10512), .A3(g10570), .ZN(g12208) );
NOR3_X4 U_g12213 ( .A1(g10453), .A2(g10516), .A3(g10572), .ZN(g12213) );
NOR3_X4 U_g12214 ( .A1(g10457), .A2(g10518), .A3(g10580), .ZN(g12214) );
NOR3_X4 U_g12215 ( .A1(g10459), .A2(g10521), .A3(g10583), .ZN(g12215) );
NOR3_X4 U_g12216 ( .A1(g10462), .A2(g10523), .A3(g10585), .ZN(g12216) );
NOR3_X4 U_g12217 ( .A1(g10465), .A2(g10526), .A3(g10588), .ZN(g12217) );
NOR3_X4 U_g12224 ( .A1(g10469), .A2(g10528), .A3(g10589), .ZN(g12224) );
NOR3_X4 U_g12231 ( .A1(g10473), .A2(g10532), .A3(g10591), .ZN(g12231) );
NOR3_X4 U_g12232 ( .A1(g10474), .A2(g10534), .A3(g10594), .ZN(g12232) );
NOR3_X4 U_g12233 ( .A1(g10477), .A2(g10537), .A3(g10596), .ZN(g12233) );
NOR3_X4 U_g12234 ( .A1(g10479), .A2(g10540), .A3(g10599), .ZN(g12234) );
NOR3_X4 U_g12245 ( .A1(g10495), .A2(g10557), .A3(g10604), .ZN(g12245) );
NOR3_X4 U_g12247 ( .A1(g10499), .A2(g10559), .A3(g10605), .ZN(g12247) );
NOR3_X4 U_g12248 ( .A1(g10508), .A2(g10567), .A3(g10612), .ZN(g12248) );
NOR3_X4 U_g12249 ( .A1(g10510), .A2(g10568), .A3(g10613), .ZN(g12249) );
NOR3_X4 U_g12250 ( .A1(g10513), .A2(g10571), .A3(g10615), .ZN(g12250) );
NOR3_X4 U_g12262 ( .A1(g10519), .A2(g10581), .A3(g10623), .ZN(g12262) );
NOR3_X4 U_g12263 ( .A1(g10524), .A2(g10586), .A3(g10627), .ZN(g12263) );
NOR3_X4 U_g12268 ( .A1(g10529), .A2(g10590), .A3(g10629), .ZN(g12268) );
NOR3_X4 U_g12269 ( .A1(g10533), .A2(g10592), .A3(g10637), .ZN(g12269) );
NOR3_X4 U_g12270 ( .A1(g10535), .A2(g10595), .A3(g10640), .ZN(g12270) );
NOR3_X4 U_g12271 ( .A1(g10538), .A2(g10597), .A3(g10642), .ZN(g12271) );
NOR3_X4 U_g12272 ( .A1(g10541), .A2(g10600), .A3(g10645), .ZN(g12272) );
NOR3_X4 U_g12288 ( .A1(g10569), .A2(g10614), .A3(g10651), .ZN(g12288) );
NOR3_X4 U_g12290 ( .A1(g10573), .A2(g10616), .A3(g10652), .ZN(g12290) );
NOR3_X4 U_g12291 ( .A1(g10582), .A2(g10624), .A3(g10659), .ZN(g12291) );
NOR3_X4 U_g12292 ( .A1(g10584), .A2(g10625), .A3(g10660), .ZN(g12292) );
NOR3_X4 U_g12293 ( .A1(g10587), .A2(g10628), .A3(g10662), .ZN(g12293) );
NOR3_X4 U_g12305 ( .A1(g10593), .A2(g10638), .A3(g10670), .ZN(g12305) );
NOR3_X4 U_g12306 ( .A1(g10598), .A2(g10643), .A3(g10674), .ZN(g12306) );
NOR3_X4 U_g12324 ( .A1(g10626), .A2(g10661), .A3(g10681), .ZN(g12324) );
NOR3_X4 U_g12326 ( .A1(g10630), .A2(g10663), .A3(g10682), .ZN(g12326) );
NOR3_X4 U_g12327 ( .A1(g10639), .A2(g10671), .A3(g10689), .ZN(g12327) );
NOR3_X4 U_g12328 ( .A1(g10641), .A2(g10672), .A3(g10690), .ZN(g12328) );
NOR3_X4 U_g12329 ( .A1(g10644), .A2(g10675), .A3(g10692), .ZN(g12329) );
NOR3_X4 U_g12339 ( .A1(g10650), .A2(g10678), .A3(g10704), .ZN(g12339) );
NOR3_X4 U_g12352 ( .A1(g10673), .A2(g10691), .A3(g10710), .ZN(g12352) );
NOR3_X4 U_g12369 ( .A1(g10680), .A2(g10707), .A3(g10724), .ZN(g12369) );
NOR3_X4 U_g12388 ( .A1(g10709), .A2(g10727), .A3(g10745), .ZN(g12388) );
NOR3_X4 U_g12418 ( .A1(g10729), .A2(g10748), .A3(g10764), .ZN(g12418) );
NOR2_X4 U_g12431 ( .A1(g8580), .A2(g10730), .ZN(g12431) );
NOR2_X4 U_g12436 ( .A1(g8587), .A2(g10749), .ZN(g12436) );
NOR2_X4 U_g12441 ( .A1(g8594), .A2(g10767), .ZN(g12441) );
NOR2_X4 U_g12446 ( .A1(g8605), .A2(g10773), .ZN(g12446) );
NOR2_X4 U_g12451 ( .A1(g499), .A2(g8983), .ZN(g12451) );
NOR3_X4 U_g12457 ( .A1(g9009), .A2(g9033), .A3(g9048), .ZN(g12457) );
NOR3_X4 U_g12467 ( .A1(g9034), .A2(g9056), .A3(g9065), .ZN(g12467) );
NOR3_X4 U_g12482 ( .A1(g9057), .A2(g9073), .A3(g9082), .ZN(g12482) );
NOR3_X4 U_g12487 ( .A1(g10108), .A2(g10198), .A3(g10283), .ZN(g12487) );
NOR3_X4 U_g12499 ( .A1(g9074), .A2(g9090), .A3(g9101), .ZN(g12499) );
NOR3_X4 U_g12507 ( .A1(g10213), .A2(g10300), .A3(g10376), .ZN(g12507) );
NOR3_X4 U_g12524 ( .A1(g10315), .A2(g10393), .A3(g10455), .ZN(g12524) );
NOR3_X4 U_g12539 ( .A1(g10408), .A2(g10472), .A3(g10531), .ZN(g12539) );
NOR3_X4 U_g12698 ( .A1(g11347), .A2(g11420), .A3(g8327), .ZN(g12698) );
NOR3_X4 U_g12747 ( .A1(g11421), .A2(g8328), .A3(g8385), .ZN(g12747) );
NOR3_X4 U_g12755 ( .A1(g11431), .A2(g8339), .A3(g8394), .ZN(g12755) );
NOR2_X4 U_g12780 ( .A1(g9187), .A2(g9161), .ZN(g12780) );
NOR3_X4 U_g12781 ( .A1(g8329), .A2(g8386), .A3(g8431), .ZN(g12781) );
NOR3_X4 U_g12789 ( .A1(g8340), .A2(g8395), .A3(g8437), .ZN(g12789) );
NOR3_X4 U_g12797 ( .A1(g8350), .A2(g8406), .A3(g8446), .ZN(g12797) );
NOR3_X4 U_g12814 ( .A1(g8387), .A2(g8432), .A3(g8463), .ZN(g12814) );
NOR2_X4 U_g12819 ( .A1(g9248), .A2(g9203), .ZN(g12819) );
NOR3_X4 U_g12820 ( .A1(g8396), .A2(g8438), .A3(g8466), .ZN(g12820) );
NOR3_X4 U_g12828 ( .A1(g8407), .A2(g8447), .A3(g8472), .ZN(g12828) );
NOR3_X4 U_g12836 ( .A1(g8417), .A2(g8458), .A3(g8481), .ZN(g12836) );
NOR3_X4 U_g12849 ( .A1(g8433), .A2(g8464), .A3(g8485), .ZN(g12849) );
NOR3_X4 U_g12852 ( .A1(g8439), .A2(g8467), .A3(g8488), .ZN(g12852) );
NOR2_X4 U_g12857 ( .A1(g9326), .A2(g9264), .ZN(g12857) );
NOR3_X4 U_g12858 ( .A1(g8448), .A2(g8473), .A3(g8491), .ZN(g12858) );
NOR3_X4 U_g12866 ( .A1(g8459), .A2(g8482), .A3(g8497), .ZN(g12866) );
NOR3_X4 U_g12880 ( .A1(g8465), .A2(g8486), .A3(g8502), .ZN(g12880) );
NOR2_X4 U_g12883 ( .A1(g10038), .A2(g6284), .ZN(g12883) );
NOR3_X4 U_g12890 ( .A1(g8468), .A2(g8489), .A3(g8505), .ZN(g12890) );
NOR3_X4 U_g12893 ( .A1(g8474), .A2(g8492), .A3(g8508), .ZN(g12893) );
NOR2_X4 U_g12898 ( .A1(g9407), .A2(g9342), .ZN(g12898) );
NOR3_X4 U_g12899 ( .A1(g8483), .A2(g8498), .A3(g8511), .ZN(g12899) );
NOR3_X4 U_g12912 ( .A1(g8484), .A2(g8500), .A3(g8515), .ZN(g12912) );
NOR3_X4 U_g12913 ( .A1(g8487), .A2(g8503), .A3(g8518), .ZN(g12913) );
NOR3_X4 U_g12920 ( .A1(g8490), .A2(g8506), .A3(g8521), .ZN(g12920) );
NOR2_X4 U_g12923 ( .A1(g10147), .A2(g6421), .ZN(g12923) );
NOR3_X4 U_g12930 ( .A1(g8493), .A2(g8509), .A3(g8524), .ZN(g12930) );
NOR3_X4 U_g12933 ( .A1(g8499), .A2(g8512), .A3(g8527), .ZN(g12933) );
NOR3_X4 U_g12939 ( .A1(g8501), .A2(g8516), .A3(g8531), .ZN(g12939) );
NOR3_X4 U_g12941 ( .A1(g8504), .A2(g8519), .A3(g8534), .ZN(g12941) );
NOR3_X4 U_g12942 ( .A1(g8507), .A2(g8522), .A3(g8537), .ZN(g12942) );
NOR3_X4 U_g12949 ( .A1(g8510), .A2(g8525), .A3(g8540), .ZN(g12949) );
NOR2_X4 U_g12952 ( .A1(g10252), .A2(g6626), .ZN(g12952) );
NOR3_X4 U_g12959 ( .A1(g8513), .A2(g8528), .A3(g8543), .ZN(g12959) );
NOR3_X4 U_g12967 ( .A1(g8517), .A2(g8532), .A3(g8546), .ZN(g12967) );
NOR3_X4 U_g12968 ( .A1(g8520), .A2(g8535), .A3(g8548), .ZN(g12968) );
NOR3_X4 U_g12970 ( .A1(g8523), .A2(g8538), .A3(g8551), .ZN(g12970) );
NOR3_X4 U_g12971 ( .A1(g8526), .A2(g8541), .A3(g8554), .ZN(g12971) );
NOR3_X4 U_g12978 ( .A1(g8529), .A2(g8544), .A3(g8557), .ZN(g12978) );
NOR2_X4 U_g12981 ( .A1(g10354), .A2(g6890), .ZN(g12981) );
NOR3_X4 U_g12991 ( .A1(g8536), .A2(g8549), .A3(g8559), .ZN(g12991) );
NOR3_X4 U_g12992 ( .A1(g8539), .A2(g8552), .A3(g8561), .ZN(g12992) );
NOR3_X4 U_g12994 ( .A1(g8542), .A2(g8555), .A3(g8564), .ZN(g12994) );
NOR3_X4 U_g12995 ( .A1(g8545), .A2(g8558), .A3(g8567), .ZN(g12995) );
NOR3_X4 U_g13001 ( .A1(g8553), .A2(g8562), .A3(g8570), .ZN(g13001) );
NOR3_X4 U_g13002 ( .A1(g8556), .A2(g8565), .A3(g8572), .ZN(g13002) );
NOR3_X4 U_g13022 ( .A1(g8566), .A2(g8573), .A3(g8576), .ZN(g13022) );
NOR4_X4 U_g13024 ( .A1(g11481), .A2(g8045), .A3(g7928), .A4(g7880), .ZN(g13024) );
NOR3_X4 U_g13111 ( .A1(g8601), .A2(g8612), .A3(g8621), .ZN(g13111) );
NOR3_X4 U_g13124 ( .A1(g8613), .A2(g8625), .A3(g8631), .ZN(g13124) );
NOR3_X4 U_g13135 ( .A1(g8626), .A2(g8635), .A3(g8650), .ZN(g13135) );
NOR3_X4 U_g13143 ( .A1(g8636), .A2(g8654), .A3(g8666), .ZN(g13143) );
NOR3_X4 U_g13149 ( .A1(g8676), .A2(g8687), .A3(g8703), .ZN(g13149) );
NOR3_X4 U_g13155 ( .A1(g8688), .A2(g8705), .A3(g8722), .ZN(g13155) );
NOR3_X4 U_g13160 ( .A1(g8704), .A2(g8717), .A3(g8751), .ZN(g13160) );
NOR3_X4 U_g13164 ( .A1(g8706), .A2(g8724), .A3(g8760), .ZN(g13164) );
NOR3_X4 U_g13171 ( .A1(g8723), .A2(g8755), .A3(g8774), .ZN(g13171) );
NOR3_X4 U_g13175 ( .A1(g8725), .A2(g8762), .A3(g8783), .ZN(g13175) );
NOR3_X4 U_g13182 ( .A1(g8761), .A2(g8778), .A3(g8797), .ZN(g13182) );
NOR3_X4 U_g13194 ( .A1(g8784), .A2(g8801), .A3(g8816), .ZN(g13194) );
NOR3_X4 U_g13228 ( .A1(g8841), .A2(g8861), .A3(g8892), .ZN(g13228) );
NOR3_X4 U_g13251 ( .A1(g8868), .A2(g8899), .A3(g8932), .ZN(g13251) );
NOR3_X4 U_g13274 ( .A1(g8906), .A2(g8939), .A3(g8972), .ZN(g13274) );
NOR4_X4 U_g13286 ( .A1(g11481), .A2(g11332), .A3(g11190), .A4(g7880), .ZN(g13286) );
NOR3_X4 U_g13299 ( .A1(g8946), .A2(g8979), .A3(g9004), .ZN(g13299) );
NOR4_X4 U_g13310 ( .A1(g11481), .A2(g11332), .A3(g11190), .A4(g11069), .ZN(g13310) );
NOR4_X4 U_g13313 ( .A1(g8183), .A2(g11332), .A3(g11190), .A4(g7880), .ZN(g13313) );
NOR4_X4 U_g13331 ( .A1(g8183), .A2(g11332), .A3(g11190), .A4(g11069), .ZN(g13331) );
NOR4_X4 U_g13332 ( .A1(g11481), .A2(g8045), .A3(g11190), .A4(g7880), .ZN(g13332) );
NOR4_X4 U_g13353 ( .A1(g11481), .A2(g8045), .A3(g11190), .A4(g11069), .ZN(g13353) );
NOR4_X4 U_g13354 ( .A1(g8183), .A2(g8045), .A3(g11190), .A4(g7880), .ZN(g13354) );
NOR4_X4 U_g13374 ( .A1(g8183), .A2(g8045), .A3(g11190), .A4(g11069), .ZN(g13374) );
NOR4_X4 U_g13375 ( .A1(g11481), .A2(g11332), .A3(g7928), .A4(g7880), .ZN(g13375) );
NOR3_X4 U_g13378 ( .A1(g9026), .A2(g9047), .A3(g9061), .ZN(g13378) );
NOR4_X4 U_g13401 ( .A1(g11481), .A2(g11332), .A3(g7928), .A4(g11069), .ZN(g13401) );
NOR4_X4 U_g13404 ( .A1(g8183), .A2(g11332), .A3(g7928), .A4(g7880), .ZN(g13404) );
NOR2_X4 U_g15661 ( .A1(g11737), .A2(g7345), .ZN(g15661) );
NOR2_X4 U_g15797 ( .A1(g13305), .A2(g7143), .ZN(g15797) );
NOR2_X4 U_g15873 ( .A1(g11617), .A2(g7562), .ZN(g15873) );
NOR2_X4 U_g15959 ( .A1(g2814), .A2(g13082), .ZN(g15959) );
NOR2_X4 U_g15978 ( .A1(g11737), .A2(g7152), .ZN(g15978) );
NOR3_X4 U_g16020 ( .A1(g6200), .A2(g12457), .A3(g10952), .ZN(g16020) );
NOR3_X4 U_g16036 ( .A1(g6289), .A2(g12467), .A3(g10952), .ZN(g16036) );
NOR3_X4 U_g16058 ( .A1(g6426), .A2(g12482), .A3(g10952), .ZN(g16058) );
NOR3_X4 U_g16082 ( .A1(g10952), .A2(g6140), .A3(g12487), .ZN(g16082) );
NOR3_X4 U_g16094 ( .A1(g6631), .A2(g12499), .A3(g10952), .ZN(g16094) );
NOR3_X4 U_g16120 ( .A1(g10952), .A2(g6161), .A3(g12507), .ZN(g16120) );
NOR3_X4 U_g16171 ( .A1(g10952), .A2(g6188), .A3(g12524), .ZN(g16171) );
NOR3_X4 U_g16230 ( .A1(g10952), .A2(g6220), .A3(g12539), .ZN(g16230) );
NOR2_X4 U_g16498 ( .A1(g14158), .A2(g14347), .ZN(g16498) );
NOR2_X4 U_g16520 ( .A1(g14273), .A2(g14459), .ZN(g16520) );
NOR2_X4 U_g16551 ( .A1(g14395), .A2(g14546), .ZN(g16551) );
NOR3_X4 U_g16567 ( .A1(g15904), .A2(g15880), .A3(g15859), .ZN(g16567) );
NOR3_X4 U_g16570 ( .A1(g15904), .A2(g15880), .A3(g14630), .ZN(g16570) );
NOR2_X4 U_g16583 ( .A1(g14507), .A2(g14601), .ZN(g16583) );
NOR3_X4 U_g16591 ( .A1(g15933), .A2(g15913), .A3(g15890), .ZN(g16591) );
NOR3_X4 U_g16594 ( .A1(g15933), .A2(g15913), .A3(g14650), .ZN(g16594) );
NOR3_X4 U_g16611 ( .A1(g15962), .A2(g15942), .A3(g15923), .ZN(g16611) );
NOR3_X4 U_g16614 ( .A1(g15962), .A2(g15942), .A3(g14677), .ZN(g16614) );
NOR3_X4 U_g16629 ( .A1(g15981), .A2(g15971), .A3(g15952), .ZN(g16629) );
NOR3_X4 U_g16632 ( .A1(g15981), .A2(g15971), .A3(g14711), .ZN(g16632) );
NOR3_X4 U_g16643 ( .A1(g15904), .A2(g14642), .A3(g15859), .ZN(g16643) );
NOR2_X4 U_g16654 ( .A1(g14690), .A2(g12477), .ZN(g16654) );
NOR3_X4 U_g16655 ( .A1(g15933), .A2(g14669), .A3(g15890), .ZN(g16655) );
NOR2_X4 U_g16671 ( .A1(g14724), .A2(g12494), .ZN(g16671) );
NOR3_X4 U_g16672 ( .A1(g15962), .A2(g14703), .A3(g15923), .ZN(g16672) );
NOR2_X4 U_g16679 ( .A1(g14797), .A2(g14895), .ZN(g16679) );
NOR2_X4 U_g16692 ( .A1(g14752), .A2(g12514), .ZN(g16692) );
NOR3_X4 U_g16693 ( .A1(g15981), .A2(g14737), .A3(g15952), .ZN(g16693) );
NOR2_X4 U_g16705 ( .A1(g14849), .A2(g14976), .ZN(g16705) );
NOR2_X4 U_g16718 ( .A1(g14773), .A2(g12531), .ZN(g16718) );
NOR2_X4 U_g16736 ( .A1(g14922), .A2(g15065), .ZN(g16736) );
NOR2_X4 U_g16778 ( .A1(g15003), .A2(g15161), .ZN(g16778) );
NOR2_X4 U_g16802 ( .A1(g13469), .A2(g3897), .ZN(g16802) );
NOR2_X4 U_g16803 ( .A1(g15593), .A2(g12908), .ZN(g16803) );
NOR2_X4 U_g16823 ( .A1(g5362), .A2(g13469), .ZN(g16823) );
NOR2_X4 U_g16824 ( .A1(g15658), .A2(g12938), .ZN(g16824) );
NOR2_X4 U_g16829 ( .A1(g14956), .A2(g12564), .ZN(g16829) );
NOR2_X4 U_g16835 ( .A1(g15717), .A2(g12966), .ZN(g16835) );
NOR2_X4 U_g16841 ( .A1(g15021), .A2(g12607), .ZN(g16841) );
NOR2_X4 U_g16844 ( .A1(g15754), .A2(g12989), .ZN(g16844) );
NOR2_X4 U_g16845 ( .A1(g15755), .A2(g12990), .ZN(g16845) );
NOR2_X4 U_g16847 ( .A1(g15095), .A2(g12650), .ZN(g16847) );
NOR2_X4 U_g16851 ( .A1(g15781), .A2(g13000), .ZN(g16851) );
NOR2_X4 U_g16853 ( .A1(g15801), .A2(g13009), .ZN(g16853) );
NOR2_X4 U_g16854 ( .A1(g15802), .A2(g13010), .ZN(g16854) );
NOR2_X4 U_g16857 ( .A1(g15817), .A2(g13023), .ZN(g16857) );
NOR2_X4 U_g16860 ( .A1(g15828), .A2(g13031), .ZN(g16860) );
NOR2_X4 U_g16861 ( .A1(g15829), .A2(g13032), .ZN(g16861) );
NOR2_X4 U_g16866 ( .A1(g15840), .A2(g13042), .ZN(g16866) );
NOR2_X4 U_g16880 ( .A1(g15852), .A2(g13056), .ZN(g16880) );
NOR3_X4 U_g17012 ( .A1(g14657), .A2(g14642), .A3(g15859), .ZN(g17012) );
NOR3_X4 U_g17025 ( .A1(g15904), .A2(g15880), .A3(g15859), .ZN(g17025) );
NOR3_X4 U_g17042 ( .A1(g14691), .A2(g14669), .A3(g15890), .ZN(g17042) );
NOR3_X4 U_g17051 ( .A1(g14657), .A2(g15880), .A3(g14630), .ZN(g17051) );
NOR3_X4 U_g17059 ( .A1(g15933), .A2(g15913), .A3(g15890), .ZN(g17059) );
NOR3_X4 U_g17076 ( .A1(g14725), .A2(g14703), .A3(g15923), .ZN(g17076) );
NOR3_X4 U_g17086 ( .A1(g14691), .A2(g15913), .A3(g14650), .ZN(g17086) );
NOR3_X4 U_g17094 ( .A1(g15962), .A2(g15942), .A3(g15923), .ZN(g17094) );
NOR3_X4 U_g17111 ( .A1(g14753), .A2(g14737), .A3(g15952), .ZN(g17111) );
NOR3_X4 U_g17124 ( .A1(g14725), .A2(g15942), .A3(g14677), .ZN(g17124) );
NOR3_X4 U_g17132 ( .A1(g15981), .A2(g15971), .A3(g15952), .ZN(g17132) );
NOR3_X4 U_g17151 ( .A1(g14753), .A2(g15971), .A3(g14711), .ZN(g17151) );
NOR2_X4 U_g17186 ( .A1(g7949), .A2(g14144), .ZN(g17186) );
NOR2_X4 U_g17197 ( .A1(g8000), .A2(g14259), .ZN(g17197) );
NOR2_X4 U_g17204 ( .A1(g8075), .A2(g14381), .ZN(g17204) );
NOR2_X4 U_g17209 ( .A1(g8160), .A2(g14493), .ZN(g17209) );
NOR2_X4 U_g17213 ( .A1(g4326), .A2(g14442), .ZN(g17213) );
NOR2_X4 U_g17215 ( .A1(g15904), .A2(g14642), .ZN(g17215) );
NOR2_X4 U_g17216 ( .A1(g4495), .A2(g14529), .ZN(g17216) );
NOR2_X4 U_g17218 ( .A1(g15933), .A2(g14669), .ZN(g17218) );
NOR2_X4 U_g17219 ( .A1(g4671), .A2(g14584), .ZN(g17219) );
NOR2_X4 U_g17220 ( .A1(g15962), .A2(g14703), .ZN(g17220) );
NOR2_X4 U_g17221 ( .A1(g4848), .A2(g14618), .ZN(g17221) );
NOR2_X4 U_g17222 ( .A1(g15998), .A2(g16003), .ZN(g17222) );
NOR2_X4 U_g17223 ( .A1(g15981), .A2(g14737), .ZN(g17223) );
NOR2_X4 U_g17224 ( .A1(g16004), .A2(g16009), .ZN(g17224) );
NOR2_X4 U_g17225 ( .A1(g16008), .A2(g16015), .ZN(g17225) );
NOR2_X4 U_g17226 ( .A1(g16010), .A2(g16017), .ZN(g17226) );
NOR2_X4 U_g17228 ( .A1(g16016), .A2(g16029), .ZN(g17228) );
NOR2_X4 U_g17229 ( .A1(g16019), .A2(g16032), .ZN(g17229) );
NOR2_X4 U_g17234 ( .A1(g16028), .A2(g16045), .ZN(g17234) );
NOR2_X4 U_g17235 ( .A1(g16030), .A2(g16047), .ZN(g17235) );
NOR2_X4 U_g17236 ( .A1(g16033), .A2(g16051), .ZN(g17236) );
NOR2_X4 U_g17246 ( .A1(g16046), .A2(g16066), .ZN(g17246) );
NOR2_X4 U_g17247 ( .A1(g16050), .A2(g16070), .ZN(g17247) );
NOR2_X4 U_g17248 ( .A1(g16052), .A2(g16072), .ZN(g17248) );
NOR2_X4 U_g17269 ( .A1(g16067), .A2(g16100), .ZN(g17269) );
NOR2_X4 U_g17270 ( .A1(g16071), .A2(g16104), .ZN(g17270) );
NOR2_X4 U_g17271 ( .A1(g16073), .A2(g16106), .ZN(g17271) );
NOR2_X4 U_g17302 ( .A1(g16103), .A2(g16135), .ZN(g17302) );
NOR2_X4 U_g17303 ( .A1(g16105), .A2(g16137), .ZN(g17303) );
NOR2_X4 U_g17340 ( .A1(g16136), .A2(g16183), .ZN(g17340) );
NOR2_X4 U_g17341 ( .A1(g16138), .A2(g16185), .ZN(g17341) );
NOR2_X4 U_g17383 ( .A1(g16184), .A2(g16238), .ZN(g17383) );
NOR2_X4 U_g17429 ( .A1(g16239), .A2(g16288), .ZN(g17429) );
NOR2_X4 U_g17507 ( .A1(g16298), .A2(g13318), .ZN(g17507) );
NOR2_X4 U_g17896 ( .A1(g14352), .A2(g16020), .ZN(g17896) );
NOR2_X4 U_g18007 ( .A1(g14464), .A2(g16036), .ZN(g18007) );
NOR2_X4 U_g18085 ( .A1(g16085), .A2(g6363), .ZN(g18085) );
NOR2_X4 U_g18124 ( .A1(g14551), .A2(g16058), .ZN(g18124) );
NOR2_X4 U_g18201 ( .A1(g16123), .A2(g6568), .ZN(g18201) );
NOR2_X4 U_g18240 ( .A1(g14606), .A2(g16094), .ZN(g18240) );
NOR2_X4 U_g18308 ( .A1(g16174), .A2(g6832), .ZN(g18308) );
NOR2_X4 U_g18352 ( .A1(g16082), .A2(g14249), .ZN(g18352) );
NOR2_X4 U_g18401 ( .A1(g16233), .A2(g7134), .ZN(g18401) );
NOR2_X4 U_g18430 ( .A1(g16020), .A2(g14352), .ZN(g18430) );
NOR2_X4 U_g18447 ( .A1(g16120), .A2(g14371), .ZN(g18447) );
NOR2_X4 U_g18503 ( .A1(g16036), .A2(g14464), .ZN(g18503) );
NOR2_X4 U_g18520 ( .A1(g16171), .A2(g14483), .ZN(g18520) );
NOR2_X4 U_g18548 ( .A1(g14249), .A2(g16082), .ZN(g18548) );
NOR2_X4 U_g18567 ( .A1(g16058), .A2(g14551), .ZN(g18567) );
NOR2_X4 U_g18584 ( .A1(g16230), .A2(g14570), .ZN(g18584) );
NOR2_X4 U_g18590 ( .A1(g16439), .A2(g7522), .ZN(g18590) );
NOR2_X4 U_g18598 ( .A1(g14371), .A2(g16120), .ZN(g18598) );
NOR2_X4 U_g18617 ( .A1(g16094), .A2(g14606), .ZN(g18617) );
NOR2_X4 U_g18623 ( .A1(g15902), .A2(g2814), .ZN(g18623) );
NOR2_X4 U_g18626 ( .A1(g16463), .A2(g7549), .ZN(g18626) );
NOR2_X4 U_g18630 ( .A1(g14483), .A2(g16171), .ZN(g18630) );
NOR2_X4 U_g18639 ( .A1(g14570), .A2(g16230), .ZN(g18639) );
NOR2_X4 U_g18669 ( .A1(g13623), .A2(g13634), .ZN(g18669) );
NOR2_X4 U_g18678 ( .A1(g13625), .A2(g11771), .ZN(g18678) );
NOR2_X4 U_g18707 ( .A1(g13636), .A2(g11788), .ZN(g18707) );
NOR2_X4 U_g18719 ( .A1(g13643), .A2(g13656), .ZN(g18719) );
NOR2_X4 U_g18726 ( .A1(g13645), .A2(g11805), .ZN(g18726) );
NOR2_X4 U_g18743 ( .A1(g13648), .A2(g11814), .ZN(g18743) );
NOR2_X4 U_g18754 ( .A1(g13655), .A2(g11816), .ZN(g18754) );
NOR2_X4 U_g18755 ( .A1(g13871), .A2(g12274), .ZN(g18755) );
NOR2_X4 U_g18763 ( .A1(g13671), .A2(g11838), .ZN(g18763) );
NOR2_X4 U_g18780 ( .A1(g13674), .A2(g11847), .ZN(g18780) );
NOR2_X4 U_g18781 ( .A1(g13675), .A2(g11851), .ZN(g18781) );
NOR2_X4 U_g18782 ( .A1(g13676), .A2(g13705), .ZN(g18782) );
NOR2_X4 U_g18794 ( .A1(g13701), .A2(g11880), .ZN(g18794) );
NOR2_X4 U_g18803 ( .A1(g13704), .A2(g11885), .ZN(g18803) );
NOR2_X4 U_g18804 ( .A1(g13905), .A2(g12331), .ZN(g18804) );
NOR2_X4 U_g18820 ( .A1(g13738), .A2(g11922), .ZN(g18820) );
NOR2_X4 U_g18821 ( .A1(g13740), .A2(g11926), .ZN(g18821) );
NOR2_X4 U_g18835 ( .A1(g13788), .A2(g11966), .ZN(g18835) );
NOR2_X4 U_g18836 ( .A1(g13789), .A2(g11967), .ZN(g18836) );
NOR2_X4 U_g18837 ( .A1(g13998), .A2(g12376), .ZN(g18837) );
NOR2_X4 U_g18852 ( .A1(g13815), .A2(g12012), .ZN(g18852) );
NOR2_X4 U_g18866 ( .A1(g13834), .A2(g12069), .ZN(g18866) );
NOR2_X4 U_g18867 ( .A1(g13835), .A2(g12070), .ZN(g18867) );
NOR2_X4 U_g18868 ( .A1(g14143), .A2(g12419), .ZN(g18868) );
NOR2_X4 U_g18883 ( .A1(g13846), .A2(g12128), .ZN(g18883) );
NOR2_X4 U_g18885 ( .A1(g13847), .A2(g12129), .ZN(g18885) );
NOR2_X4 U_g18906 ( .A1(g13855), .A2(g12186), .ZN(g18906) );
NOR2_X4 U_g18907 ( .A1(g14336), .A2(g12429), .ZN(g18907) );
NOR2_X4 U_g18942 ( .A1(g13870), .A2(g12273), .ZN(g18942) );
NOR2_X4 U_g18957 ( .A1(g13884), .A2(g12307), .ZN(g18957) );
NOR2_X4 U_g18968 ( .A1(g13904), .A2(g12330), .ZN(g18968) );
NOR2_X4 U_g18975 ( .A1(g13944), .A2(g12353), .ZN(g18975) );
NOR2_X4 U_g19144 ( .A1(g17268), .A2(g14884), .ZN(g19144) );
NOR2_X4 U_g19149 ( .A1(g17339), .A2(g15020), .ZN(g19149) );
NOR2_X4 U_g19153 ( .A1(g17381), .A2(g15093), .ZN(g19153) );
NOR2_X4 U_g19154 ( .A1(g17382), .A2(g15094), .ZN(g19154) );
NOR2_X4 U_g19157 ( .A1(g17428), .A2(g15171), .ZN(g19157) );
NOR2_X4 U_g19160 ( .A1(g17446), .A2(g15178), .ZN(g19160) );
NOR2_X4 U_g19162 ( .A1(g17485), .A2(g15243), .ZN(g19162) );
NOR2_X4 U_g19163 ( .A1(g17486), .A2(g15244), .ZN(g19163) );
NOR2_X4 U_g19165 ( .A1(g17526), .A2(g15264), .ZN(g19165) );
NOR2_X4 U_g19167 ( .A1(g17556), .A2(g15320), .ZN(g19167) );
NOR2_X4 U_g19171 ( .A1(g17616), .A2(g15356), .ZN(g19171) );
NOR2_X4 U_g19172 ( .A1(g17635), .A2(g15388), .ZN(g19172) );
NOR2_X4 U_g19173 ( .A1(g17636), .A2(g15389), .ZN(g19173) );
NOR2_X4 U_g19177 ( .A1(g17713), .A2(g15442), .ZN(g19177) );
NOR2_X4 U_g19178 ( .A1(g17718), .A2(g15452), .ZN(g19178) );
NOR2_X4 U_g19179 ( .A1(g17719), .A2(g15453), .ZN(g19179) );
NOR2_X4 U_g19184 ( .A1(g17798), .A2(g15520), .ZN(g19184) );
NOR2_X4 U_g19219 ( .A1(g18165), .A2(g15753), .ZN(g19219) );
NOR2_X4 U_g20008 ( .A1(g18977), .A2(g7338), .ZN(g20008) );
NOR2_X4 U_g20054 ( .A1(g19001), .A2(g16867), .ZN(g20054) );
NOR2_X4 U_g20095 ( .A1(g16507), .A2(g16895), .ZN(g20095) );
NOR2_X4 U_g20120 ( .A1(g16529), .A2(g16924), .ZN(g20120) );
NOR2_X4 U_g20150 ( .A1(g16560), .A2(g16954), .ZN(g20150) );
NOR2_X4 U_g20153 ( .A1(g16536), .A2(g7583), .ZN(g20153) );
NOR2_X4 U_g20299 ( .A1(g16665), .A2(g16884), .ZN(g20299) );
NOR2_X4 U_g20310 ( .A1(g16850), .A2(g13654), .ZN(g20310) );
NOR2_X4 U_g20314 ( .A1(g13646), .A2(g16855), .ZN(g20314) );
NOR2_X4 U_g20318 ( .A1(g16686), .A2(g16913), .ZN(g20318) );
NOR2_X4 U_g20333 ( .A1(g13672), .A2(g16859), .ZN(g20333) );
NOR2_X4 U_g20337 ( .A1(g16712), .A2(g16943), .ZN(g20337) );
NOR2_X4 U_g20343 ( .A1(g16856), .A2(g13703), .ZN(g20343) );
NOR2_X4 U_g20353 ( .A1(g13702), .A2(g16864), .ZN(g20353) );
NOR2_X4 U_g20357 ( .A1(g16743), .A2(g16974), .ZN(g20357) );
NOR2_X4 U_g20375 ( .A1(g13739), .A2(g16879), .ZN(g20375) );
NOR2_X4 U_g20376 ( .A1(g16865), .A2(g13787), .ZN(g20376) );
NOR2_X4 U_g20417 ( .A1(g16907), .A2(g13833), .ZN(g20417) );
NOR2_X4 U_g20682 ( .A1(g19160), .A2(g10024), .ZN(g20682) );
NOR2_X4 U_g20717 ( .A1(g19165), .A2(g10133), .ZN(g20717) );
NOR2_X4 U_g20752 ( .A1(g19171), .A2(g10238), .ZN(g20752) );
NOR2_X4 U_g20789 ( .A1(g19177), .A2(g10340), .ZN(g20789) );
NOR2_X4 U_g20841 ( .A1(g14767), .A2(g19552), .ZN(g20841) );
NOR2_X4 U_g20874 ( .A1(g17301), .A2(g19594), .ZN(g20874) );
NOR2_X4 U_g20875 ( .A1(g19584), .A2(g17352), .ZN(g20875) );
NOR2_X4 U_g20876 ( .A1(g19585), .A2(g17353), .ZN(g20876) );
NOR2_X4 U_g20877 ( .A1(g3919), .A2(g19830), .ZN(g20877) );
NOR2_X4 U_g20878 ( .A1(g19600), .A2(g17395), .ZN(g20878) );
NOR2_X4 U_g20879 ( .A1(g19601), .A2(g17396), .ZN(g20879) );
NOR2_X4 U_g20880 ( .A1(g19602), .A2(g17397), .ZN(g20880) );
NOR2_X4 U_g20881 ( .A1(g19603), .A2(g17398), .ZN(g20881) );
NOR2_X4 U_g20882 ( .A1(g19614), .A2(g17408), .ZN(g20882) );
NOR2_X4 U_g20883 ( .A1(g19615), .A2(g17409), .ZN(g20883) );
NOR2_X4 U_g20884 ( .A1(g5394), .A2(g19830), .ZN(g20884) );
NOR2_X4 U_g20891 ( .A1(g19626), .A2(g17447), .ZN(g20891) );
NOR2_X4 U_g20892 ( .A1(g19627), .A2(g17448), .ZN(g20892) );
NOR2_X4 U_g20893 ( .A1(g19628), .A2(g17449), .ZN(g20893) );
NOR2_X4 U_g20894 ( .A1(g19629), .A2(g17450), .ZN(g20894) );
NOR2_X4 U_g20895 ( .A1(g19633), .A2(g17461), .ZN(g20895) );
NOR2_X4 U_g20896 ( .A1(g19634), .A2(g17462), .ZN(g20896) );
NOR2_X4 U_g20897 ( .A1(g19635), .A2(g17463), .ZN(g20897) );
NOR2_X4 U_g20898 ( .A1(g19636), .A2(g17464), .ZN(g20898) );
NOR2_X4 U_g20899 ( .A1(g19647), .A2(g17474), .ZN(g20899) );
NOR2_X4 U_g20900 ( .A1(g19648), .A2(g17475), .ZN(g20900) );
NOR2_X4 U_g20901 ( .A1(g19660), .A2(g17508), .ZN(g20901) );
NOR2_X4 U_g20902 ( .A1(g19661), .A2(g17509), .ZN(g20902) );
NOR2_X4 U_g20903 ( .A1(g19662), .A2(g17510), .ZN(g20903) );
NOR2_X4 U_g20910 ( .A1(g19666), .A2(g17527), .ZN(g20910) );
NOR2_X4 U_g20911 ( .A1(g19667), .A2(g17528), .ZN(g20911) );
NOR2_X4 U_g20912 ( .A1(g19668), .A2(g17529), .ZN(g20912) );
NOR2_X4 U_g20913 ( .A1(g19669), .A2(g17530), .ZN(g20913) );
NOR2_X4 U_g20914 ( .A1(g19673), .A2(g17541), .ZN(g20914) );
NOR2_X4 U_g20915 ( .A1(g19674), .A2(g17542), .ZN(g20915) );
NOR2_X4 U_g20916 ( .A1(g19675), .A2(g17543), .ZN(g20916) );
NOR2_X4 U_g20917 ( .A1(g19676), .A2(g17544), .ZN(g20917) );
NOR2_X4 U_g20918 ( .A1(g19687), .A2(g17554), .ZN(g20918) );
NOR2_X4 U_g20919 ( .A1(g19688), .A2(g17555), .ZN(g20919) );
NOR2_X4 U_g20920 ( .A1(g19691), .A2(g19726), .ZN(g20920) );
NOR2_X4 U_g20921 ( .A1(g19697), .A2(g17576), .ZN(g20921) );
NOR2_X4 U_g20922 ( .A1(g19698), .A2(g17577), .ZN(g20922) );
NOR2_X4 U_g20923 ( .A1(g19699), .A2(g17578), .ZN(g20923) );
NOR2_X4 U_g20924 ( .A1(g19700), .A2(g15257), .ZN(g20924) );
NOR2_X4 U_g20925 ( .A1(g19708), .A2(g17598), .ZN(g20925) );
NOR2_X4 U_g20926 ( .A1(g19709), .A2(g17599), .ZN(g20926) );
NOR2_X4 U_g20927 ( .A1(g19710), .A2(g17600), .ZN(g20927) );
NOR2_X4 U_g20934 ( .A1(g19714), .A2(g17617), .ZN(g20934) );
NOR2_X4 U_g20935 ( .A1(g19715), .A2(g17618), .ZN(g20935) );
NOR2_X4 U_g20936 ( .A1(g19716), .A2(g17619), .ZN(g20936) );
NOR2_X4 U_g20937 ( .A1(g19717), .A2(g17620), .ZN(g20937) );
NOR2_X4 U_g20938 ( .A1(g19721), .A2(g17631), .ZN(g20938) );
NOR2_X4 U_g20939 ( .A1(g19722), .A2(g17632), .ZN(g20939) );
NOR2_X4 U_g20940 ( .A1(g19723), .A2(g17633), .ZN(g20940) );
NOR2_X4 U_g20941 ( .A1(g19724), .A2(g17634), .ZN(g20941) );
NOR2_X4 U_g20944 ( .A1(g19731), .A2(g17652), .ZN(g20944) );
NOR2_X4 U_g20945 ( .A1(g19732), .A2(g17653), .ZN(g20945) );
NOR2_X4 U_g20946 ( .A1(g19733), .A2(g17654), .ZN(g20946) );
NOR2_X4 U_g20947 ( .A1(g19734), .A2(g15335), .ZN(g20947) );
NOR2_X4 U_g20948 ( .A1(g19735), .A2(g15336), .ZN(g20948) );
NOR2_X4 U_g20949 ( .A1(g19741), .A2(g17673), .ZN(g20949) );
NOR2_X4 U_g20950 ( .A1(g19742), .A2(g17674), .ZN(g20950) );
NOR2_X4 U_g20951 ( .A1(g19743), .A2(g17675), .ZN(g20951) );
NOR2_X4 U_g20952 ( .A1(g19744), .A2(g15349), .ZN(g20952) );
NOR2_X4 U_g20953 ( .A1(g19752), .A2(g17695), .ZN(g20953) );
NOR2_X4 U_g20954 ( .A1(g19753), .A2(g17696), .ZN(g20954) );
NOR2_X4 U_g20955 ( .A1(g19754), .A2(g17697), .ZN(g20955) );
NOR2_X4 U_g20962 ( .A1(g19758), .A2(g17714), .ZN(g20962) );
NOR2_X4 U_g20963 ( .A1(g19759), .A2(g17715), .ZN(g20963) );
NOR2_X4 U_g20964 ( .A1(g19760), .A2(g17716), .ZN(g20964) );
NOR2_X4 U_g20965 ( .A1(g19761), .A2(g17717), .ZN(g20965) );
NOR2_X4 U_g20966 ( .A1(g19765), .A2(g17734), .ZN(g20966) );
NOR2_X4 U_g20967 ( .A1(g19766), .A2(g17735), .ZN(g20967) );
NOR2_X4 U_g20968 ( .A1(g19767), .A2(g17736), .ZN(g20968) );
NOR2_X4 U_g20969 ( .A1(g19768), .A2(g15402), .ZN(g20969) );
NOR2_X4 U_g20970 ( .A1(g19769), .A2(g15403), .ZN(g20970) );
NOR2_X4 U_g20972 ( .A1(g19774), .A2(g17752), .ZN(g20972) );
NOR2_X4 U_g20973 ( .A1(g19775), .A2(g17753), .ZN(g20973) );
NOR2_X4 U_g20974 ( .A1(g19776), .A2(g17754), .ZN(g20974) );
NOR2_X4 U_g20975 ( .A1(g19777), .A2(g15421), .ZN(g20975) );
NOR2_X4 U_g20976 ( .A1(g19778), .A2(g15422), .ZN(g20976) );
NOR2_X4 U_g20977 ( .A1(g19784), .A2(g17773), .ZN(g20977) );
NOR2_X4 U_g20978 ( .A1(g19785), .A2(g17774), .ZN(g20978) );
NOR2_X4 U_g20979 ( .A1(g19786), .A2(g17775), .ZN(g20979) );
NOR2_X4 U_g20980 ( .A1(g19787), .A2(g15435), .ZN(g20980) );
NOR2_X4 U_g20981 ( .A1(g19795), .A2(g17795), .ZN(g20981) );
NOR2_X4 U_g20982 ( .A1(g19796), .A2(g17796), .ZN(g20982) );
NOR2_X4 U_g20983 ( .A1(g19797), .A2(g17797), .ZN(g20983) );
NOR2_X4 U_g20989 ( .A1(g19802), .A2(g17812), .ZN(g20989) );
NOR2_X4 U_g20990 ( .A1(g19803), .A2(g17813), .ZN(g20990) );
NOR2_X4 U_g20991 ( .A1(g19804), .A2(g17814), .ZN(g20991) );
NOR2_X4 U_g20992 ( .A1(g19805), .A2(g15470), .ZN(g20992) );
NOR2_X4 U_g20993 ( .A1(g19807), .A2(g17835), .ZN(g20993) );
NOR2_X4 U_g20994 ( .A1(g19808), .A2(g17836), .ZN(g20994) );
NOR2_X4 U_g20995 ( .A1(g19809), .A2(g17837), .ZN(g20995) );
NOR2_X4 U_g20996 ( .A1(g19810), .A2(g15486), .ZN(g20996) );
NOR2_X4 U_g20997 ( .A1(g19811), .A2(g15487), .ZN(g20997) );
NOR2_X4 U_g20999 ( .A1(g19816), .A2(g17853), .ZN(g20999) );
NOR2_X4 U_g21000 ( .A1(g19817), .A2(g17854), .ZN(g21000) );
NOR2_X4 U_g21001 ( .A1(g19818), .A2(g17855), .ZN(g21001) );
NOR2_X4 U_g21002 ( .A1(g19819), .A2(g15505), .ZN(g21002) );
NOR2_X4 U_g21003 ( .A1(g19820), .A2(g15506), .ZN(g21003) );
NOR2_X4 U_g21004 ( .A1(g19826), .A2(g17874), .ZN(g21004) );
NOR2_X4 U_g21005 ( .A1(g19827), .A2(g17875), .ZN(g21005) );
NOR2_X4 U_g21006 ( .A1(g19828), .A2(g17876), .ZN(g21006) );
NOR2_X4 U_g21007 ( .A1(g19829), .A2(g15519), .ZN(g21007) );
NOR2_X4 U_g21008 ( .A1(g19836), .A2(g17877), .ZN(g21008) );
NOR2_X4 U_g21009 ( .A1(g19839), .A2(g17900), .ZN(g21009) );
NOR2_X4 U_g21010 ( .A1(g19840), .A2(g17901), .ZN(g21010) );
NOR2_X4 U_g21011 ( .A1(g19841), .A2(g17902), .ZN(g21011) );
NOR2_X4 U_g21015 ( .A1(g19846), .A2(g17924), .ZN(g21015) );
NOR2_X4 U_g21016 ( .A1(g19847), .A2(g17925), .ZN(g21016) );
NOR2_X4 U_g21017 ( .A1(g19848), .A2(g17926), .ZN(g21017) );
NOR2_X4 U_g21018 ( .A1(g19849), .A2(g15556), .ZN(g21018) );
NOR2_X4 U_g21019 ( .A1(g19851), .A2(g17947), .ZN(g21019) );
NOR2_X4 U_g21020 ( .A1(g19852), .A2(g17948), .ZN(g21020) );
NOR2_X4 U_g21021 ( .A1(g19853), .A2(g17949), .ZN(g21021) );
NOR2_X4 U_g21022 ( .A1(g19854), .A2(g15572), .ZN(g21022) );
NOR2_X4 U_g21023 ( .A1(g19855), .A2(g15573), .ZN(g21023) );
NOR2_X4 U_g21025 ( .A1(g19860), .A2(g17965), .ZN(g21025) );
NOR2_X4 U_g21026 ( .A1(g19861), .A2(g17966), .ZN(g21026) );
NOR2_X4 U_g21027 ( .A1(g19862), .A2(g17967), .ZN(g21027) );
NOR2_X4 U_g21028 ( .A1(g19863), .A2(g15591), .ZN(g21028) );
NOR2_X4 U_g21029 ( .A1(g19864), .A2(g15592), .ZN(g21029) );
NOR2_X4 U_g21031 ( .A1(g19869), .A2(g17989), .ZN(g21031) );
NOR2_X4 U_g21032 ( .A1(g19870), .A2(g17990), .ZN(g21032) );
NOR2_X4 U_g21033 ( .A1(g19872), .A2(g18011), .ZN(g21033) );
NOR2_X4 U_g21034 ( .A1(g19873), .A2(g18012), .ZN(g21034) );
NOR2_X4 U_g21035 ( .A1(g19874), .A2(g18013), .ZN(g21035) );
NOR2_X4 U_g21039 ( .A1(g19879), .A2(g18035), .ZN(g21039) );
NOR2_X4 U_g21040 ( .A1(g19880), .A2(g18036), .ZN(g21040) );
NOR2_X4 U_g21041 ( .A1(g19881), .A2(g18037), .ZN(g21041) );
NOR2_X4 U_g21042 ( .A1(g19882), .A2(g15634), .ZN(g21042) );
NOR2_X4 U_g21043 ( .A1(g19884), .A2(g18058), .ZN(g21043) );
NOR2_X4 U_g21044 ( .A1(g19885), .A2(g18059), .ZN(g21044) );
NOR2_X4 U_g21045 ( .A1(g19886), .A2(g18060), .ZN(g21045) );
NOR2_X4 U_g21046 ( .A1(g19887), .A2(g15650), .ZN(g21046) );
NOR2_X4 U_g21047 ( .A1(g19888), .A2(g15651), .ZN(g21047) );
NOR2_X4 U_g21048 ( .A1(g19889), .A2(g18062), .ZN(g21048) );
NOR2_X4 U_g21051 ( .A1(g19895), .A2(g18088), .ZN(g21051) );
NOR2_X4 U_g21052 ( .A1(g19900), .A2(g18106), .ZN(g21052) );
NOR2_X4 U_g21053 ( .A1(g19901), .A2(g18107), .ZN(g21053) );
NOR2_X4 U_g21054 ( .A1(g19903), .A2(g18128), .ZN(g21054) );
NOR2_X4 U_g21055 ( .A1(g19904), .A2(g18129), .ZN(g21055) );
NOR2_X4 U_g21056 ( .A1(g19905), .A2(g18130), .ZN(g21056) );
NOR2_X4 U_g21060 ( .A1(g19910), .A2(g18152), .ZN(g21060) );
NOR2_X4 U_g21061 ( .A1(g19911), .A2(g18153), .ZN(g21061) );
NOR2_X4 U_g21062 ( .A1(g19912), .A2(g18154), .ZN(g21062) );
NOR2_X4 U_g21063 ( .A1(g19913), .A2(g15710), .ZN(g21063) );
NOR2_X4 U_g21065 ( .A1(g19914), .A2(g18169), .ZN(g21065) );
NOR2_X4 U_g21070 ( .A1(g19920), .A2(g18204), .ZN(g21070) );
NOR2_X4 U_g21071 ( .A1(g19925), .A2(g18222), .ZN(g21071) );
NOR2_X4 U_g21072 ( .A1(g19926), .A2(g18223), .ZN(g21072) );
NOR2_X4 U_g21073 ( .A1(g19928), .A2(g18244), .ZN(g21073) );
NOR2_X4 U_g21074 ( .A1(g19929), .A2(g18245), .ZN(g21074) );
NOR2_X4 U_g21075 ( .A1(g19930), .A2(g18246), .ZN(g21075) );
NOR2_X4 U_g21080 ( .A1(g19935), .A2(g18311), .ZN(g21080) );
NOR2_X4 U_g21081 ( .A1(g19940), .A2(g18329), .ZN(g21081) );
NOR2_X4 U_g21082 ( .A1(g19941), .A2(g18330), .ZN(g21082) );
NOR2_X4 U_g21083 ( .A1(g19943), .A2(g18333), .ZN(g21083) );
NOR2_X4 U_g21084 ( .A1(g20011), .A2(g20048), .ZN(g21084) );
NOR2_X4 U_g21094 ( .A1(g19952), .A2(g18404), .ZN(g21094) );
NOR3_X4 U_g21095 ( .A1(g20012), .A2(g20049), .A3(g20084), .ZN(g21095) );
NOR3_X4 U_g21096 ( .A1(g20013), .A2(g20051), .A3(g20087), .ZN(g21096) );
NOR3_X4 U_g21104 ( .A1(g20050), .A2(g20085), .A3(g20106), .ZN(g21104) );
NOR3_X4 U_g21105 ( .A1(g20052), .A2(g20088), .A3(g20109), .ZN(g21105) );
NOR3_X4 U_g21106 ( .A1(g20053), .A2(g20090), .A3(g20112), .ZN(g21106) );
NOR3_X4 U_g21116 ( .A1(g20086), .A2(g20107), .A3(g20131), .ZN(g21116) );
NOR3_X4 U_g21117 ( .A1(g20089), .A2(g20110), .A3(g20133), .ZN(g21117) );
NOR3_X4 U_g21118 ( .A1(g20091), .A2(g20113), .A3(g20136), .ZN(g21118) );
NOR3_X4 U_g21119 ( .A1(g20092), .A2(g20115), .A3(g20139), .ZN(g21119) );
NOR3_X4 U_g21133 ( .A1(g20108), .A2(g20132), .A3(g20156), .ZN(g21133) );
NOR3_X4 U_g21134 ( .A1(g20111), .A2(g20134), .A3(g20157), .ZN(g21134) );
NOR3_X4 U_g21135 ( .A1(g20114), .A2(g20137), .A3(g20160), .ZN(g21135) );
NOR3_X4 U_g21147 ( .A1(g20135), .A2(g20158), .A3(g20188), .ZN(g21147) );
NOR3_X4 U_g21148 ( .A1(g20138), .A2(g20161), .A3(g20190), .ZN(g21148) );
NOR2_X4 U_g21149 ( .A1(g20015), .A2(g19981), .ZN(g21149) );
NOR2_X4 U_g21167 ( .A1(g20159), .A2(g20189), .ZN(g21167) );
NOR3_X4 U_g21168 ( .A1(g20162), .A2(g20191), .A3(g20220), .ZN(g21168) );
NOR2_X4 U_g21169 ( .A1(g20057), .A2(g20019), .ZN(g21169) );
NOR2_X4 U_g21183 ( .A1(g20192), .A2(g20221), .ZN(g21183) );
NOR2_X4 U_g21189 ( .A1(g20098), .A2(g20061), .ZN(g21189) );
NOR2_X4 U_g21204 ( .A1(g20123), .A2(g20102), .ZN(g21204) );
NOR2_X4 U_g21211 ( .A1(g19240), .A2(g19230), .ZN(g21211) );
NOR2_X4 U_g21219 ( .A1(g19253), .A2(g19243), .ZN(g21219) );
NOR3_X4 U_g21227 ( .A1(g18414), .A2(g18485), .A3(g20295), .ZN(g21227) );
NOR2_X4 U_g21228 ( .A1(g19388), .A2(g17118), .ZN(g21228) );
NOR2_X4 U_g21230 ( .A1(g19266), .A2(g19256), .ZN(g21230) );
NOR2_X4 U_g21233 ( .A1(g19418), .A2(g17145), .ZN(g21233) );
NOR2_X4 U_g21235 ( .A1(g19281), .A2(g19269), .ZN(g21235) );
NOR2_X4 U_g21238 ( .A1(g19954), .A2(g5890), .ZN(g21238) );
NOR2_X4 U_g21242 ( .A1(g19455), .A2(g17168), .ZN(g21242) );
NOR2_X4 U_g21246 ( .A1(g19984), .A2(g5929), .ZN(g21246) );
NOR2_X4 U_g21250 ( .A1(g19482), .A2(g17183), .ZN(g21250) );
NOR2_X4 U_g21255 ( .A1(g20022), .A2(g5963), .ZN(g21255) );
NOR2_X4 U_g21263 ( .A1(g20064), .A2(g5992), .ZN(g21263) );
NOR2_X4 U_g21316 ( .A1(g20460), .A2(g16111), .ZN(g21316) );
NOR2_X4 U_g21331 ( .A1(g20472), .A2(g16153), .ZN(g21331) );
NOR2_X4 U_g21346 ( .A1(g20480), .A2(g13247), .ZN(g21346) );
NOR2_X4 U_g21364 ( .A1(g20486), .A2(g13266), .ZN(g21364) );
NOR2_X4 U_g21385 ( .A1(g20492), .A2(g13289), .ZN(g21385) );
NOR2_X4 U_g21407 ( .A1(g20499), .A2(g13316), .ZN(g21407) );
NOR2_X4 U_g21432 ( .A1(g20502), .A2(g13335), .ZN(g21432) );
NOR2_X4 U_g21435 ( .A1(g20503), .A2(g16385), .ZN(g21435) );
NOR2_X4 U_g21467 ( .A1(g20506), .A2(g13355), .ZN(g21467) );
NOR2_X4 U_g21470 ( .A1(g20512), .A2(g16417), .ZN(g21470) );
NOR2_X4 U_g21502 ( .A1(g20525), .A2(g16445), .ZN(g21502) );
NOR2_X4 U_g21615 ( .A1(g16567), .A2(g19957), .ZN(g21615) );
NOR3_X4 U_g21618 ( .A1(g20016), .A2(g14079), .A3(g14165), .ZN(g21618) );
NOR2_X4 U_g21636 ( .A1(g20473), .A2(g6513), .ZN(g21636) );
NOR2_X4 U_g21643 ( .A1(g16591), .A2(g19987), .ZN(g21643) );
NOR3_X4 U_g21646 ( .A1(g20058), .A2(g14194), .A3(g14280), .ZN(g21646) );
NOR2_X4 U_g21665 ( .A1(g20507), .A2(g18352), .ZN(g21665) );
NOR2_X4 U_g21667 ( .A1(g20481), .A2(g6777), .ZN(g21667) );
NOR2_X4 U_g21674 ( .A1(g16611), .A2(g20025), .ZN(g21674) );
NOR3_X4 U_g21677 ( .A1(g20099), .A2(g14309), .A3(g14402), .ZN(g21677) );
NOR2_X4 U_g21694 ( .A1(g20526), .A2(g18447), .ZN(g21694) );
NOR2_X4 U_g21696 ( .A1(g20487), .A2(g7079), .ZN(g21696) );
NOR2_X4 U_g21703 ( .A1(g16629), .A2(g20067), .ZN(g21703) );
NOR3_X4 U_g21706 ( .A1(g20124), .A2(g14431), .A3(g14514), .ZN(g21706) );
NOR2_X4 U_g21711 ( .A1(g19830), .A2(g15780), .ZN(g21711) );
NOR2_X4 U_g21730 ( .A1(g20545), .A2(g18520), .ZN(g21730) );
NOR2_X4 U_g21732 ( .A1(g20493), .A2(g7329), .ZN(g21732) );
NOR3_X4 U_g21738 ( .A1(g19444), .A2(g17893), .A3(g14079), .ZN(g21738) );
NOR2_X4 U_g21739 ( .A1(g20507), .A2(g18430), .ZN(g21739) );
NOR2_X4 U_g21756 ( .A1(g19070), .A2(g18584), .ZN(g21756) );
NOR3_X4 U_g21762 ( .A1(g19471), .A2(g18004), .A3(g14194), .ZN(g21762) );
NOR2_X4 U_g21763 ( .A1(g20526), .A2(g18503), .ZN(g21763) );
NOR3_X4 U_g21778 ( .A1(g19494), .A2(g18121), .A3(g14309), .ZN(g21778) );
NOR2_X4 U_g21779 ( .A1(g20545), .A2(g18567), .ZN(g21779) );
NOR3_X4 U_g21793 ( .A1(g19515), .A2(g18237), .A3(g14431), .ZN(g21793) );
NOR2_X4 U_g21794 ( .A1(g19070), .A2(g18617), .ZN(g21794) );
NOR2_X4 U_g21796 ( .A1(g19830), .A2(g13004), .ZN(g21796) );
NOR2_X4 U_g21842 ( .A1(g13609), .A2(g19150), .ZN(g21842) );
NOR2_X4 U_g21843 ( .A1(g13619), .A2(g19155), .ZN(g21843) );
NOR2_X4 U_g21845 ( .A1(g13631), .A2(g19161), .ZN(g21845) );
NOR2_X4 U_g21847 ( .A1(g13642), .A2(g19166), .ZN(g21847) );
NOR2_X4 U_g21851 ( .A1(g19252), .A2(g8842), .ZN(g21851) );
NOR2_X4 U_g21878 ( .A1(g16964), .A2(g19228), .ZN(g21878) );
NOR2_X4 U_g21880 ( .A1(g13854), .A2(g19236), .ZN(g21880) );
NOR2_X4 U_g21882 ( .A1(g13862), .A2(g19248), .ZN(g21882) );
NOR2_X4 U_g21884 ( .A1(g19260), .A2(g19284), .ZN(g21884) );
NOR2_X4 U_g21887 ( .A1(g13519), .A2(g19289), .ZN(g21887) );
NOR2_X4 U_g21889 ( .A1(g19285), .A2(g19316), .ZN(g21889) );
NOR2_X4 U_g21890 ( .A1(g13530), .A2(g19307), .ZN(g21890) );
NOR2_X4 U_g21893 ( .A1(g13541), .A2(g19328), .ZN(g21893) );
NOR2_X4 U_g21894 ( .A1(g19317), .A2(g19356), .ZN(g21894) );
NOR2_X4 U_g21901 ( .A1(g13552), .A2(g19355), .ZN(g21901) );
NOR2_X4 U_g21968 ( .A1(g21234), .A2(g19476), .ZN(g21968) );
NOR2_X4 U_g21969 ( .A1(g20895), .A2(g10133), .ZN(g21969) );
NOR2_X4 U_g21970 ( .A1(g17182), .A2(g21226), .ZN(g21970) );
NOR2_X4 U_g21971 ( .A1(g21243), .A2(g19499), .ZN(g21971) );
NOR2_X4 U_g21972 ( .A1(g20914), .A2(g10238), .ZN(g21972) );
NOR2_X4 U_g21973 ( .A1(g21251), .A2(g19520), .ZN(g21973) );
NOR2_X4 U_g21974 ( .A1(g20938), .A2(g10340), .ZN(g21974) );
NOR2_X4 U_g21975 ( .A1(g21245), .A2(g21259), .ZN(g21975) );
NOR3_X4 U_g21980 ( .A1(g21252), .A2(g19531), .A3(g19540), .ZN(g21980) );
NOR2_X4 U_g21981 ( .A1(g21254), .A2(g21267), .ZN(g21981) );
NOR3_X4 U_g21987 ( .A1(g21260), .A2(g19541), .A3(g19544), .ZN(g21987) );
NOR2_X4 U_g21988 ( .A1(g21262), .A2(g21276), .ZN(g21988) );
NOR3_X4 U_g22000 ( .A1(g21268), .A2(g19545), .A3(g19547), .ZN(g22000) );
NOR2_X4 U_g22001 ( .A1(g21270), .A2(g21283), .ZN(g22001) );
NOR3_X4 U_g22013 ( .A1(g21277), .A2(g19548), .A3(g19551), .ZN(g22013) );
NOR2_X4 U_g22025 ( .A1(g21284), .A2(g19549), .ZN(g22025) );
NOR2_X4 U_g22026 ( .A1(g21083), .A2(g18407), .ZN(g22026) );
NOR2_X4 U_g22027 ( .A1(g21290), .A2(g19553), .ZN(g22027) );
NOR2_X4 U_g22028 ( .A1(g21291), .A2(g19554), .ZN(g22028) );
NOR2_X4 U_g22029 ( .A1(g21292), .A2(g19555), .ZN(g22029) );
NOR2_X4 U_g22030 ( .A1(g21298), .A2(g19557), .ZN(g22030) );
NOR2_X4 U_g22031 ( .A1(g21299), .A2(g19558), .ZN(g22031) );
NOR2_X4 U_g22032 ( .A1(g21300), .A2(g19559), .ZN(g22032) );
NOR2_X4 U_g22033 ( .A1(g21301), .A2(g19560), .ZN(g22033) );
NOR2_X4 U_g22034 ( .A1(g21302), .A2(g19561), .ZN(g22034) );
NOR2_X4 U_g22035 ( .A1(g21303), .A2(g19562), .ZN(g22035) );
NOR2_X4 U_g22037 ( .A1(g21304), .A2(g19564), .ZN(g22037) );
NOR2_X4 U_g22038 ( .A1(g21305), .A2(g19565), .ZN(g22038) );
NOR2_X4 U_g22039 ( .A1(g21306), .A2(g19566), .ZN(g22039) );
NOR2_X4 U_g22040 ( .A1(g21307), .A2(g19567), .ZN(g22040) );
NOR2_X4 U_g22041 ( .A1(g21308), .A2(g19568), .ZN(g22041) );
NOR2_X4 U_g22042 ( .A1(g21309), .A2(g19569), .ZN(g22042) );
NOR2_X4 U_g22043 ( .A1(g21310), .A2(g19570), .ZN(g22043) );
NOR2_X4 U_g22044 ( .A1(g21311), .A2(g19571), .ZN(g22044) );
NOR2_X4 U_g22045 ( .A1(g21312), .A2(g19572), .ZN(g22045) );
NOR2_X4 U_g22047 ( .A1(g21313), .A2(g19574), .ZN(g22047) );
NOR2_X4 U_g22048 ( .A1(g21314), .A2(g19575), .ZN(g22048) );
NOR2_X4 U_g22049 ( .A1(g21315), .A2(g19576), .ZN(g22049) );
NOR2_X4 U_g22054 ( .A1(g21319), .A2(g19586), .ZN(g22054) );
NOR2_X4 U_g22055 ( .A1(g21320), .A2(g19587), .ZN(g22055) );
NOR2_X4 U_g22056 ( .A1(g21321), .A2(g19588), .ZN(g22056) );
NOR2_X4 U_g22057 ( .A1(g21322), .A2(g19589), .ZN(g22057) );
NOR2_X4 U_g22058 ( .A1(g21323), .A2(g19590), .ZN(g22058) );
NOR2_X4 U_g22059 ( .A1(g21324), .A2(g19591), .ZN(g22059) );
NOR2_X4 U_g22060 ( .A1(g21325), .A2(g19592), .ZN(g22060) );
NOR2_X4 U_g22061 ( .A1(g21326), .A2(g19593), .ZN(g22061) );
NOR2_X4 U_g22063 ( .A1(g21328), .A2(g19597), .ZN(g22063) );
NOR2_X4 U_g22064 ( .A1(g21329), .A2(g19598), .ZN(g22064) );
NOR2_X4 U_g22065 ( .A1(g21330), .A2(g19599), .ZN(g22065) );
NOR2_X4 U_g22066 ( .A1(g21334), .A2(g19604), .ZN(g22066) );
NOR2_X4 U_g22067 ( .A1(g21335), .A2(g19605), .ZN(g22067) );
NOR2_X4 U_g22068 ( .A1(g21336), .A2(g19606), .ZN(g22068) );
NOR2_X4 U_g22073 ( .A1(g21337), .A2(g19616), .ZN(g22073) );
NOR2_X4 U_g22074 ( .A1(g21338), .A2(g19617), .ZN(g22074) );
NOR2_X4 U_g22075 ( .A1(g21339), .A2(g19618), .ZN(g22075) );
NOR2_X4 U_g22076 ( .A1(g21340), .A2(g19619), .ZN(g22076) );
NOR2_X4 U_g22077 ( .A1(g21341), .A2(g19620), .ZN(g22077) );
NOR2_X4 U_g22078 ( .A1(g21342), .A2(g19621), .ZN(g22078) );
NOR2_X4 U_g22079 ( .A1(g21343), .A2(g19623), .ZN(g22079) );
NOR2_X4 U_g22080 ( .A1(g21344), .A2(g19624), .ZN(g22080) );
NOR2_X4 U_g22081 ( .A1(g21345), .A2(g19625), .ZN(g22081) );
NOR2_X4 U_g22087 ( .A1(g21349), .A2(g19630), .ZN(g22087) );
NOR2_X4 U_g22088 ( .A1(g21350), .A2(g19631), .ZN(g22088) );
NOR2_X4 U_g22089 ( .A1(g21351), .A2(g19632), .ZN(g22089) );
NOR2_X4 U_g22090 ( .A1(g21352), .A2(g19637), .ZN(g22090) );
NOR2_X4 U_g22091 ( .A1(g21353), .A2(g19638), .ZN(g22091) );
NOR2_X4 U_g22092 ( .A1(g21354), .A2(g19639), .ZN(g22092) );
NOR2_X4 U_g22097 ( .A1(g21355), .A2(g19649), .ZN(g22097) );
NOR2_X4 U_g22098 ( .A1(g21356), .A2(g19650), .ZN(g22098) );
NOR2_X4 U_g22099 ( .A1(g21357), .A2(g19651), .ZN(g22099) );
NOR2_X4 U_g22100 ( .A1(g21360), .A2(g19653), .ZN(g22100) );
NOR2_X4 U_g22101 ( .A1(g21361), .A2(g19654), .ZN(g22101) );
NOR2_X4 U_g22102 ( .A1(g21362), .A2(g19655), .ZN(g22102) );
NOR2_X4 U_g22103 ( .A1(g21363), .A2(g19656), .ZN(g22103) );
NOR2_X4 U_g22104 ( .A1(g21367), .A2(g19663), .ZN(g22104) );
NOR2_X4 U_g22105 ( .A1(g21368), .A2(g19664), .ZN(g22105) );
NOR2_X4 U_g22106 ( .A1(g21369), .A2(g19665), .ZN(g22106) );
NOR2_X4 U_g22112 ( .A1(g21370), .A2(g19670), .ZN(g22112) );
NOR2_X4 U_g22113 ( .A1(g21371), .A2(g19671), .ZN(g22113) );
NOR2_X4 U_g22114 ( .A1(g21372), .A2(g19672), .ZN(g22114) );
NOR2_X4 U_g22115 ( .A1(g21373), .A2(g19677), .ZN(g22115) );
NOR2_X4 U_g22116 ( .A1(g21374), .A2(g19678), .ZN(g22116) );
NOR2_X4 U_g22117 ( .A1(g21375), .A2(g19679), .ZN(g22117) );
NOR2_X4 U_g22122 ( .A1(g21378), .A2(g19692), .ZN(g22122) );
NOR2_X4 U_g22123 ( .A1(g21379), .A2(g19693), .ZN(g22123) );
NOR2_X4 U_g22124 ( .A1(g21380), .A2(g19694), .ZN(g22124) );
NOR2_X4 U_g22125 ( .A1(g21381), .A2(g19695), .ZN(g22125) );
NOR2_X4 U_g22126 ( .A1(g21389), .A2(g19701), .ZN(g22126) );
NOR2_X4 U_g22127 ( .A1(g21390), .A2(g19702), .ZN(g22127) );
NOR2_X4 U_g22128 ( .A1(g21391), .A2(g19703), .ZN(g22128) );
NOR2_X4 U_g22129 ( .A1(g21392), .A2(g19704), .ZN(g22129) );
NOR2_X4 U_g22130 ( .A1(g21393), .A2(g19711), .ZN(g22130) );
NOR2_X4 U_g22131 ( .A1(g21394), .A2(g19712), .ZN(g22131) );
NOR2_X4 U_g22132 ( .A1(g21395), .A2(g19713), .ZN(g22132) );
NOR2_X4 U_g22138 ( .A1(g21396), .A2(g19718), .ZN(g22138) );
NOR2_X4 U_g22139 ( .A1(g21397), .A2(g19719), .ZN(g22139) );
NOR2_X4 U_g22140 ( .A1(g21398), .A2(g19720), .ZN(g22140) );
NOR2_X4 U_g22141 ( .A1(g21401), .A2(g19727), .ZN(g22141) );
NOR2_X4 U_g22142 ( .A1(g21402), .A2(g19728), .ZN(g22142) );
NOR2_X4 U_g22143 ( .A1(g21403), .A2(g19729), .ZN(g22143) );
NOR2_X4 U_g22144 ( .A1(g21410), .A2(g19730), .ZN(g22144) );
NOR2_X4 U_g22145 ( .A1(g21411), .A2(g19736), .ZN(g22145) );
NOR2_X4 U_g22146 ( .A1(g21412), .A2(g19737), .ZN(g22146) );
NOR2_X4 U_g22147 ( .A1(g21413), .A2(g19738), .ZN(g22147) );
NOR2_X4 U_g22148 ( .A1(g21414), .A2(g19739), .ZN(g22148) );
NOR2_X4 U_g22149 ( .A1(g21419), .A2(g19745), .ZN(g22149) );
NOR2_X4 U_g22150 ( .A1(g21420), .A2(g19746), .ZN(g22150) );
NOR2_X4 U_g22151 ( .A1(g21421), .A2(g19747), .ZN(g22151) );
NOR2_X4 U_g22152 ( .A1(g21422), .A2(g19748), .ZN(g22152) );
NOR2_X4 U_g22153 ( .A1(g21423), .A2(g19755), .ZN(g22153) );
NOR2_X4 U_g22154 ( .A1(g21424), .A2(g19756), .ZN(g22154) );
NOR2_X4 U_g22155 ( .A1(g21425), .A2(g19757), .ZN(g22155) );
NOR2_X4 U_g22161 ( .A1(g21428), .A2(g19764), .ZN(g22161) );
NOR2_X4 U_g22162 ( .A1(g21438), .A2(g19770), .ZN(g22162) );
NOR2_X4 U_g22163 ( .A1(g21439), .A2(g19771), .ZN(g22163) );
NOR2_X4 U_g22164 ( .A1(g21440), .A2(g19772), .ZN(g22164) );
NOR2_X4 U_g22165 ( .A1(g21444), .A2(g19773), .ZN(g22165) );
NOR2_X4 U_g22166 ( .A1(g21445), .A2(g19779), .ZN(g22166) );
NOR2_X4 U_g22167 ( .A1(g21446), .A2(g19780), .ZN(g22167) );
NOR2_X4 U_g22168 ( .A1(g21447), .A2(g19781), .ZN(g22168) );
NOR2_X4 U_g22169 ( .A1(g21448), .A2(g19782), .ZN(g22169) );
NOR2_X4 U_g22170 ( .A1(g21453), .A2(g19788), .ZN(g22170) );
NOR2_X4 U_g22171 ( .A1(g21454), .A2(g19789), .ZN(g22171) );
NOR2_X4 U_g22172 ( .A1(g21455), .A2(g19790), .ZN(g22172) );
NOR2_X4 U_g22173 ( .A1(g21456), .A2(g19791), .ZN(g22173) );
NOR2_X4 U_g22174 ( .A1(g19868), .A2(g21593), .ZN(g22174) );
NOR2_X4 U_g22177 ( .A1(g21476), .A2(g19806), .ZN(g22177) );
NOR2_X4 U_g22178 ( .A1(g21480), .A2(g19812), .ZN(g22178) );
NOR2_X4 U_g22179 ( .A1(g21481), .A2(g19813), .ZN(g22179) );
NOR2_X4 U_g22180 ( .A1(g21482), .A2(g19814), .ZN(g22180) );
NOR2_X4 U_g22181 ( .A1(g21486), .A2(g19815), .ZN(g22181) );
NOR2_X4 U_g22182 ( .A1(g21487), .A2(g19821), .ZN(g22182) );
NOR2_X4 U_g22183 ( .A1(g21488), .A2(g19822), .ZN(g22183) );
NOR2_X4 U_g22184 ( .A1(g21489), .A2(g19823), .ZN(g22184) );
NOR2_X4 U_g22185 ( .A1(g21490), .A2(g19824), .ZN(g22185) );
NOR2_X4 U_g22186 ( .A1(g21497), .A2(g19837), .ZN(g22186) );
NOR2_X4 U_g22189 ( .A1(g19899), .A2(g21622), .ZN(g22189) );
NOR2_X4 U_g22191 ( .A1(g21517), .A2(g19850), .ZN(g22191) );
NOR2_X4 U_g22192 ( .A1(g21521), .A2(g19856), .ZN(g22192) );
NOR2_X4 U_g22193 ( .A1(g21522), .A2(g19857), .ZN(g22193) );
NOR2_X4 U_g22194 ( .A1(g21523), .A2(g19858), .ZN(g22194) );
NOR2_X4 U_g22195 ( .A1(g21527), .A2(g19859), .ZN(g22195) );
NOR2_X4 U_g22198 ( .A1(g19924), .A2(g21650), .ZN(g22198) );
NOR2_X4 U_g22200 ( .A1(g21553), .A2(g19883), .ZN(g22200) );
NOR2_X4 U_g22204 ( .A1(g19939), .A2(g21681), .ZN(g22204) );
NOR2_X4 U_g22210 ( .A1(g21610), .A2(g19932), .ZN(g22210) );
NOR2_X4 U_g22216 ( .A1(g21635), .A2(g19944), .ZN(g22216) );
NOR2_X4 U_g22218 ( .A1(g21639), .A2(g19949), .ZN(g22218) );
NOR2_X4 U_g22227 ( .A1(g21658), .A2(g19953), .ZN(g22227) );
NOR2_X4 U_g22231 ( .A1(g21666), .A2(g19971), .ZN(g22231) );
NOR2_X4 U_g22234 ( .A1(g21670), .A2(g19976), .ZN(g22234) );
NOR2_X4 U_g22242 ( .A1(g21687), .A2(g19983), .ZN(g22242) );
NOR2_X4 U_g22247 ( .A1(g21695), .A2(g20001), .ZN(g22247) );
NOR2_X4 U_g22249 ( .A1(g21699), .A2(g20006), .ZN(g22249) );
NOR2_X4 U_g22263 ( .A1(g21723), .A2(g20021), .ZN(g22263) );
NOR2_X4 U_g22267 ( .A1(g21731), .A2(g20039), .ZN(g22267) );
NOR2_X4 U_g22269 ( .A1(g21735), .A2(g20044), .ZN(g22269) );
NOR2_X4 U_g22280 ( .A1(g21749), .A2(g20063), .ZN(g22280) );
NOR2_X4 U_g22284 ( .A1(g21757), .A2(g20081), .ZN(g22284) );
NOR2_X4 U_g22288 ( .A1(g20144), .A2(g21805), .ZN(g22288) );
NOR2_X4 U_g22299 ( .A1(g21773), .A2(g20104), .ZN(g22299) );
NOR2_X4 U_g22308 ( .A1(g20182), .A2(g21812), .ZN(g22308) );
NOR2_X4 U_g22336 ( .A1(g20216), .A2(g21818), .ZN(g22336) );
NOR2_X4 U_g22361 ( .A1(g20246), .A2(g21822), .ZN(g22361) );
NOR2_X4 U_g22454 ( .A1(g17012), .A2(g21891), .ZN(g22454) );
NOR2_X4 U_g22493 ( .A1(g17042), .A2(g21899), .ZN(g22493) );
NOR2_X4 U_g22536 ( .A1(g17076), .A2(g21911), .ZN(g22536) );
NOR2_X4 U_g22576 ( .A1(g17111), .A2(g21925), .ZN(g22576) );
NOR2_X4 U_g22578 ( .A1(g21892), .A2(g18982), .ZN(g22578) );
NOR2_X4 U_g22615 ( .A1(g21900), .A2(g18990), .ZN(g22615) );
NOR2_X4 U_g22651 ( .A1(g21912), .A2(g18997), .ZN(g22651) );
NOR2_X4 U_g22687 ( .A1(g21926), .A2(g19010), .ZN(g22687) );
NOR2_X4 U_g22755 ( .A1(g21271), .A2(g20842), .ZN(g22755) );
NOR2_X4 U_g22784 ( .A1(g16075), .A2(g20885), .ZN(g22784) );
NOR2_X4 U_g22789 ( .A1(g21278), .A2(g20850), .ZN(g22789) );
NOR3_X4 U_g22810 ( .A1(g16075), .A2(g20842), .A3(g21271), .ZN(g22810) );
NOR2_X4 U_g22826 ( .A1(g16113), .A2(g20904), .ZN(g22826) );
NOR2_X4 U_g22831 ( .A1(g21285), .A2(g20858), .ZN(g22831) );
NOR3_X4 U_g22851 ( .A1(g16113), .A2(g20850), .A3(g21278), .ZN(g22851) );
NOR2_X4 U_g22865 ( .A1(g16164), .A2(g20928), .ZN(g22865) );
NOR2_X4 U_g22870 ( .A1(g21293), .A2(g20866), .ZN(g22870) );
NOR3_X4 U_g22886 ( .A1(g16164), .A2(g20858), .A3(g21285), .ZN(g22886) );
NOR2_X4 U_g22900 ( .A1(g16223), .A2(g20956), .ZN(g22900) );
NOR3_X4 U_g22921 ( .A1(g16223), .A2(g20866), .A3(g21293), .ZN(g22921) );
NOR2_X4 U_g22935 ( .A1(g21903), .A2(g7466), .ZN(g22935) );
NOR2_X4 U_g22953 ( .A1(g20700), .A2(g7595), .ZN(g22953) );
NOR2_X4 U_g22985 ( .A1(g21618), .A2(g21049), .ZN(g22985) );
NOR2_X4 U_g22987 ( .A1(g21646), .A2(g21068), .ZN(g22987) );
NOR2_X4 U_g22990 ( .A1(g21677), .A2(g21078), .ZN(g22990) );
NOR2_X4 U_g22997 ( .A1(g21706), .A2(g21092), .ZN(g22997) );
NOR2_X4 U_g22999 ( .A1(g21085), .A2(g19241), .ZN(g22999) );
NOR2_X4 U_g23000 ( .A1(g16909), .A2(g21067), .ZN(g23000) );
NOR2_X4 U_g23009 ( .A1(g21738), .A2(g21107), .ZN(g23009) );
NOR2_X4 U_g23013 ( .A1(g21097), .A2(g19254), .ZN(g23013) );
NOR2_X4 U_g23014 ( .A1(g16939), .A2(g21077), .ZN(g23014) );
NOR2_X4 U_g23022 ( .A1(g16968), .A2(g21086), .ZN(g23022) );
NOR3_X4 U_g23023 ( .A1(g14256), .A2(g14175), .A3(g21123), .ZN(g23023) );
NOR2_X4 U_g23025 ( .A1(g21762), .A2(g21124), .ZN(g23025) );
NOR2_X4 U_g23029 ( .A1(g21111), .A2(g19267), .ZN(g23029) );
NOR2_X4 U_g23030 ( .A1(g16970), .A2(g21091), .ZN(g23030) );
NOR2_X4 U_g23039 ( .A1(g16989), .A2(g21098), .ZN(g23039) );
NOR3_X4 U_g23040 ( .A1(g14378), .A2(g14290), .A3(g21142), .ZN(g23040) );
NOR2_X4 U_g23042 ( .A1(g21778), .A2(g21143), .ZN(g23042) );
NOR2_X4 U_g23046 ( .A1(g21128), .A2(g19282), .ZN(g23046) );
NOR2_X4 U_g23047 ( .A1(g16991), .A2(g21103), .ZN(g23047) );
NOR2_X4 U_g23051 ( .A1(g21121), .A2(g21153), .ZN(g23051) );
NOR2_X4 U_g23058 ( .A1(g16999), .A2(g21112), .ZN(g23058) );
NOR3_X4 U_g23059 ( .A1(g14490), .A2(g14412), .A3(g21162), .ZN(g23059) );
NOR2_X4 U_g23061 ( .A1(g21793), .A2(g21163), .ZN(g23061) );
NOR3_X4 U_g23066 ( .A1(g21138), .A2(g19303), .A3(g19320), .ZN(g23066) );
NOR2_X4 U_g23067 ( .A1(g17015), .A2(g21122), .ZN(g23067) );
NOR2_X4 U_g23070 ( .A1(g21140), .A2(g21173), .ZN(g23070) );
NOR2_X4 U_g23076 ( .A1(g17023), .A2(g21129), .ZN(g23076) );
NOR3_X4 U_g23077 ( .A1(g14577), .A2(g14524), .A3(g21182), .ZN(g23077) );
NOR3_X4 U_g23080 ( .A1(g21158), .A2(g19324), .A3(g19347), .ZN(g23080) );
NOR2_X4 U_g23081 ( .A1(g17045), .A2(g21141), .ZN(g23081) );
NOR2_X4 U_g23083 ( .A1(g21160), .A2(g21193), .ZN(g23083) );
NOR2_X4 U_g23092 ( .A1(g17055), .A2(g21154), .ZN(g23092) );
NOR2_X4 U_g23093 ( .A1(g17056), .A2(g21155), .ZN(g23093) );
NOR3_X4 U_g23096 ( .A1(g21178), .A2(g19351), .A3(g19381), .ZN(g23096) );
NOR2_X4 U_g23097 ( .A1(g17079), .A2(g21161), .ZN(g23097) );
NOR2_X4 U_g23099 ( .A1(g21180), .A2(g21208), .ZN(g23099) );
NOR2_X4 U_g23110 ( .A1(g17090), .A2(g21174), .ZN(g23110) );
NOR2_X4 U_g23111 ( .A1(g17091), .A2(g21175), .ZN(g23111) );
NOR3_X4 U_g23113 ( .A1(g21198), .A2(g19385), .A3(g19413), .ZN(g23113) );
NOR2_X4 U_g23114 ( .A1(g17114), .A2(g21181), .ZN(g23114) );
NOR2_X4 U_g23117 ( .A1(g17117), .A2(g21188), .ZN(g23117) );
NOR2_X4 U_g23123 ( .A1(g17128), .A2(g21194), .ZN(g23123) );
NOR2_X4 U_g23124 ( .A1(g17129), .A2(g21195), .ZN(g23124) );
NOR2_X4 U_g23126 ( .A1(g17144), .A2(g21203), .ZN(g23126) );
NOR2_X4 U_g23132 ( .A1(g17155), .A2(g21209), .ZN(g23132) );
NOR2_X4 U_g23133 ( .A1(g17156), .A2(g21210), .ZN(g23133) );
NOR2_X4 U_g23135 ( .A1(g21229), .A2(g19449), .ZN(g23135) );
NOR2_X4 U_g23136 ( .A1(g20878), .A2(g10024), .ZN(g23136) );
NOR2_X4 U_g23137 ( .A1(g17167), .A2(g21218), .ZN(g23137) );
NOR2_X4 U_g23324 ( .A1(g22144), .A2(g10024), .ZN(g23324) );
NOR2_X4 U_g23329 ( .A1(g22165), .A2(g10133), .ZN(g23329) );
NOR2_X4 U_g23330 ( .A1(g22186), .A2(g22777), .ZN(g23330) );
NOR2_X4 U_g23339 ( .A1(g22181), .A2(g10238), .ZN(g23339) );
NOR2_X4 U_g23348 ( .A1(g22195), .A2(g10340), .ZN(g23348) );
NOR2_X4 U_g23357 ( .A1(g22210), .A2(g20127), .ZN(g23357) );
NOR2_X4 U_g23358 ( .A1(g22227), .A2(g18407), .ZN(g23358) );
NOR2_X4 U_g23359 ( .A1(g22216), .A2(g22907), .ZN(g23359) );
NOR2_X4 U_g23385 ( .A1(g17393), .A2(g22517), .ZN(g23385) );
NOR2_X4 U_g23386 ( .A1(g22483), .A2(g21388), .ZN(g23386) );
NOR2_X4 U_g23392 ( .A1(g17460), .A2(g22557), .ZN(g23392) );
NOR2_X4 U_g23393 ( .A1(g22526), .A2(g21418), .ZN(g23393) );
NOR2_X4 U_g23399 ( .A1(g17506), .A2(g22581), .ZN(g23399) );
NOR2_X4 U_g23400 ( .A1(g17540), .A2(g22597), .ZN(g23400) );
NOR2_X4 U_g23401 ( .A1(g22566), .A2(g21452), .ZN(g23401) );
NOR2_X4 U_g23406 ( .A1(g17597), .A2(g22618), .ZN(g23406) );
NOR2_X4 U_g23407 ( .A1(g17630), .A2(g22634), .ZN(g23407) );
NOR2_X4 U_g23408 ( .A1(g22606), .A2(g21494), .ZN(g23408) );
NOR2_X4 U_g23413 ( .A1(g17694), .A2(g22654), .ZN(g23413) );
NOR2_X4 U_g23418 ( .A1(g17794), .A2(g22690), .ZN(g23418) );
NOR2_X4 U_g23427 ( .A1(g22699), .A2(g21589), .ZN(g23427) );
NOR2_X4 U_g23433 ( .A1(g22726), .A2(g21611), .ZN(g23433) );
NOR2_X4 U_g23461 ( .A1(g22841), .A2(g21707), .ZN(g23461) );
NOR2_X4 U_g23477 ( .A1(g22906), .A2(g21758), .ZN(g23477) );
NOR2_X4 U_g23497 ( .A1(g22876), .A2(g5606), .ZN(g23497) );
NOR2_X4 U_g23513 ( .A1(g22911), .A2(g5631), .ZN(g23513) );
NOR2_X4 U_g23528 ( .A1(g22936), .A2(g5659), .ZN(g23528) );
NOR2_X4 U_g23539 ( .A1(g22942), .A2(g5697), .ZN(g23539) );
NOR2_X4 U_g23545 ( .A1(g22984), .A2(g20285), .ZN(g23545) );
NOR3_X4 U_g23823 ( .A1(g23009), .A2(g18490), .A3(g4456), .ZN(g23823) );
NOR3_X4 U_g23858 ( .A1(g23025), .A2(g18554), .A3(g4632), .ZN(g23858) );
NOR3_X4 U_g23892 ( .A1(g23042), .A2(g18604), .A3(g4809), .ZN(g23892) );
NOR3_X4 U_g23913 ( .A1(g23061), .A2(g18636), .A3(g4985), .ZN(g23913) );
NOR2_X4 U_g23922 ( .A1(g4456), .A2(g22985), .ZN(g23922) );
NOR3_X4 U_g23945 ( .A1(g4456), .A2(g13565), .A3(g23009), .ZN(g23945) );
NOR2_X4 U_g23950 ( .A1(g22992), .A2(g6707), .ZN(g23950) );
NOR2_X4 U_g23954 ( .A1(g4632), .A2(g22987), .ZN(g23954) );
NOR3_X4 U_g23974 ( .A1(g4632), .A2(g13573), .A3(g23025), .ZN(g23974) );
NOR2_X4 U_g23979 ( .A1(g23003), .A2(g7009), .ZN(g23979) );
NOR2_X4 U_g23983 ( .A1(g4809), .A2(g22990), .ZN(g23983) );
NOR3_X4 U_g24004 ( .A1(g4809), .A2(g13582), .A3(g23042), .ZN(g24004) );
NOR2_X4 U_g24009 ( .A1(g23017), .A2(g7259), .ZN(g24009) );
NOR2_X4 U_g24013 ( .A1(g4985), .A2(g22997), .ZN(g24013) );
NOR3_X4 U_g24038 ( .A1(g4985), .A2(g13602), .A3(g23061), .ZN(g24038) );
NOR2_X4 U_g24043 ( .A1(g23033), .A2(g7455), .ZN(g24043) );
NOR2_X4 U_g24059 ( .A1(g21990), .A2(g20809), .ZN(g24059) );
NOR2_X4 U_g24072 ( .A1(g22004), .A2(g20826), .ZN(g24072) );
NOR2_X4 U_g24083 ( .A1(g22015), .A2(g20836), .ZN(g24083) );
NOR2_X4 U_g24092 ( .A1(g22020), .A2(g20840), .ZN(g24092) );
NOR2_X4 U_g24174 ( .A1(g16894), .A2(g22206), .ZN(g24174) );
NOR2_X4 U_g24178 ( .A1(g16908), .A2(g22211), .ZN(g24178) );
NOR2_X4 U_g24179 ( .A1(g16923), .A2(g22214), .ZN(g24179) );
NOR2_X4 U_g24181 ( .A1(g16938), .A2(g22220), .ZN(g24181) );
NOR2_X4 U_g24182 ( .A1(g16953), .A2(g22223), .ZN(g24182) );
NOR2_X4 U_g24206 ( .A1(g16966), .A2(g22228), .ZN(g24206) );
NOR2_X4 U_g24207 ( .A1(g16967), .A2(g22229), .ZN(g24207) );
NOR2_X4 U_g24208 ( .A1(g16969), .A2(g22235), .ZN(g24208) );
NOR2_X4 U_g24209 ( .A1(g16984), .A2(g22238), .ZN(g24209) );
NOR2_X4 U_g24212 ( .A1(g16987), .A2(g22244), .ZN(g24212) );
NOR2_X4 U_g24213 ( .A1(g16988), .A2(g22245), .ZN(g24213) );
NOR2_X4 U_g24214 ( .A1(g16990), .A2(g22250), .ZN(g24214) );
NOR2_X4 U_g24215 ( .A1(g16993), .A2(g22254), .ZN(g24215) );
NOR2_X4 U_g24216 ( .A1(g16994), .A2(g22255), .ZN(g24216) );
NOR2_X4 U_g24218 ( .A1(g16997), .A2(g22264), .ZN(g24218) );
NOR2_X4 U_g24219 ( .A1(g16998), .A2(g22265), .ZN(g24219) );
NOR2_X4 U_g24222 ( .A1(g17017), .A2(g22272), .ZN(g24222) );
NOR2_X4 U_g24223 ( .A1(g17018), .A2(g22273), .ZN(g24223) );
NOR2_X4 U_g24225 ( .A1(g17021), .A2(g22281), .ZN(g24225) );
NOR2_X4 U_g24226 ( .A1(g17022), .A2(g22282), .ZN(g24226) );
NOR2_X4 U_g24227 ( .A1(g22270), .A2(g21137), .ZN(g24227) );
NOR2_X4 U_g24228 ( .A1(g17028), .A2(g22285), .ZN(g24228) );
NOR2_X4 U_g24230 ( .A1(g17047), .A2(g22291), .ZN(g24230) );
NOR2_X4 U_g24231 ( .A1(g17048), .A2(g22292), .ZN(g24231) );
NOR2_X4 U_g24232 ( .A1(g22637), .A2(g22665), .ZN(g24232) );
NOR2_X4 U_g24234 ( .A1(g22289), .A2(g21157), .ZN(g24234) );
NOR2_X4 U_g24235 ( .A1(g17062), .A2(g22305), .ZN(g24235) );
NOR2_X4 U_g24237 ( .A1(g17081), .A2(g22311), .ZN(g24237) );
NOR2_X4 U_g24238 ( .A1(g17082), .A2(g22312), .ZN(g24238) );
NOR2_X4 U_g24242 ( .A1(g22309), .A2(g21177), .ZN(g24242) );
NOR2_X4 U_g24243 ( .A1(g17097), .A2(g22333), .ZN(g24243) );
NOR2_X4 U_g24249 ( .A1(g22337), .A2(g21197), .ZN(g24249) );
NOR2_X4 U_g24250 ( .A1(g17135), .A2(g22358), .ZN(g24250) );
NOR2_X4 U_g24426 ( .A1(g23386), .A2(g10024), .ZN(g24426) );
NOR2_X4 U_g24428 ( .A1(g23544), .A2(g22398), .ZN(g24428) );
NOR2_X4 U_g24430 ( .A1(g23393), .A2(g10133), .ZN(g24430) );
NOR2_X4 U_g24434 ( .A1(g23401), .A2(g10238), .ZN(g24434) );
NOR2_X4 U_g24438 ( .A1(g23408), .A2(g10340), .ZN(g24438) );
NOR2_X4 U_g24445 ( .A1(g23427), .A2(g22777), .ZN(g24445) );
NOR2_X4 U_g24446 ( .A1(g23433), .A2(g22907), .ZN(g24446) );
NOR2_X4 U_g24473 ( .A1(g23461), .A2(g18407), .ZN(g24473) );
NOR2_X4 U_g24476 ( .A1(g23477), .A2(g20127), .ZN(g24476) );
NOR2_X4 U_g24479 ( .A1(g23593), .A2(g22516), .ZN(g24479) );
NOR2_X4 U_g24480 ( .A1(g23617), .A2(g23659), .ZN(g24480) );
NOR2_X4 U_g24481 ( .A1(g23618), .A2(g19696), .ZN(g24481) );
NOR2_X4 U_g24485 ( .A1(g23625), .A2(g22556), .ZN(g24485) );
NOR2_X4 U_g24486 ( .A1(g23643), .A2(g22577), .ZN(g24486) );
NOR2_X4 U_g24487 ( .A1(g23666), .A2(g23709), .ZN(g24487) );
NOR2_X4 U_g24488 ( .A1(g23667), .A2(g19740), .ZN(g24488) );
NOR2_X4 U_g24489 ( .A1(g23674), .A2(g22596), .ZN(g24489) );
NOR2_X4 U_g24490 ( .A1(g23686), .A2(g22607), .ZN(g24490) );
NOR2_X4 U_g24491 ( .A1(g15247), .A2(g23735), .ZN(g24491) );
NOR2_X4 U_g24492 ( .A1(g23689), .A2(g22610), .ZN(g24492) );
NOR2_X4 U_g24493 ( .A1(g23693), .A2(g22614), .ZN(g24493) );
NOR2_X4 U_g24494 ( .A1(g23716), .A2(g23763), .ZN(g24494) );
NOR2_X4 U_g24495 ( .A1(g23717), .A2(g19783), .ZN(g24495) );
NOR2_X4 U_g24496 ( .A1(g23724), .A2(g22633), .ZN(g24496) );
NOR2_X4 U_g24497 ( .A1(g23734), .A2(g22638), .ZN(g24497) );
NOR2_X4 U_g24498 ( .A1(g15324), .A2(g23777), .ZN(g24498) );
NOR2_X4 U_g24499 ( .A1(g15325), .A2(g23778), .ZN(g24499) );
NOR2_X4 U_g24500 ( .A1(g23740), .A2(g22643), .ZN(g24500) );
NOR2_X4 U_g24501 ( .A1(g15339), .A2(g23790), .ZN(g24501) );
NOR2_X4 U_g24502 ( .A1(g23743), .A2(g22646), .ZN(g24502) );
NOR2_X4 U_g24503 ( .A1(g23747), .A2(g22650), .ZN(g24503) );
NOR2_X4 U_g24504 ( .A1(g23770), .A2(g23818), .ZN(g24504) );
NOR2_X4 U_g24505 ( .A1(g23771), .A2(g19825), .ZN(g24505) );
NOR2_X4 U_g24506 ( .A1(g23776), .A2(g22667), .ZN(g24506) );
NOR2_X4 U_g24507 ( .A1(g15391), .A2(g23824), .ZN(g24507) );
NOR2_X4 U_g24508 ( .A1(g15392), .A2(g23825), .ZN(g24508) );
NOR2_X4 U_g24509 ( .A1(g23789), .A2(g22674), .ZN(g24509) );
NOR2_X4 U_g24510 ( .A1(g15410), .A2(g23830), .ZN(g24510) );
NOR2_X4 U_g24511 ( .A1(g15411), .A2(g23831), .ZN(g24511) );
NOR2_X4 U_g24512 ( .A1(g23795), .A2(g22679), .ZN(g24512) );
NOR2_X4 U_g24513 ( .A1(g15425), .A2(g23843), .ZN(g24513) );
NOR2_X4 U_g24514 ( .A1(g23798), .A2(g22682), .ZN(g24514) );
NOR2_X4 U_g24515 ( .A1(g23802), .A2(g22686), .ZN(g24515) );
NOR2_X4 U_g24516 ( .A1(g23820), .A2(g22700), .ZN(g24516) );
NOR2_X4 U_g24517 ( .A1(g23822), .A2(g22701), .ZN(g24517) );
NOR2_X4 U_g24519 ( .A1(g15459), .A2(g23855), .ZN(g24519) );
NOR2_X4 U_g24520 ( .A1(g23829), .A2(g22707), .ZN(g24520) );
NOR2_X4 U_g24521 ( .A1(g15475), .A2(g23859), .ZN(g24521) );
NOR2_X4 U_g24522 ( .A1(g15476), .A2(g23860), .ZN(g24522) );
NOR2_X4 U_g24523 ( .A1(g23842), .A2(g22714), .ZN(g24523) );
NOR2_X4 U_g24524 ( .A1(g15494), .A2(g23865), .ZN(g24524) );
NOR2_X4 U_g24525 ( .A1(g15495), .A2(g23866), .ZN(g24525) );
NOR2_X4 U_g24526 ( .A1(g23848), .A2(g22719), .ZN(g24526) );
NOR2_X4 U_g24527 ( .A1(g15509), .A2(g23878), .ZN(g24527) );
NOR2_X4 U_g24528 ( .A1(g23851), .A2(g22722), .ZN(g24528) );
NOR2_X4 U_g24530 ( .A1(g23857), .A2(g22732), .ZN(g24530) );
NOR2_X4 U_g24532 ( .A1(g15545), .A2(g23889), .ZN(g24532) );
NOR2_X4 U_g24533 ( .A1(g23864), .A2(g22738), .ZN(g24533) );
NOR2_X4 U_g24534 ( .A1(g15561), .A2(g23893), .ZN(g24534) );
NOR2_X4 U_g24535 ( .A1(g15562), .A2(g23894), .ZN(g24535) );
NOR2_X4 U_g24536 ( .A1(g23877), .A2(g22745), .ZN(g24536) );
NOR2_X4 U_g24537 ( .A1(g15580), .A2(g23899), .ZN(g24537) );
NOR2_X4 U_g24538 ( .A1(g15581), .A2(g23900), .ZN(g24538) );
NOR2_X4 U_g24543 ( .A1(g23891), .A2(g22764), .ZN(g24543) );
NOR2_X4 U_g24545 ( .A1(g15623), .A2(g23910), .ZN(g24545) );
NOR2_X4 U_g24546 ( .A1(g23898), .A2(g22770), .ZN(g24546) );
NOR2_X4 U_g24547 ( .A1(g15639), .A2(g23914), .ZN(g24547) );
NOR2_X4 U_g24548 ( .A1(g15640), .A2(g23915), .ZN(g24548) );
NOR2_X4 U_g24555 ( .A1(g23912), .A2(g22798), .ZN(g24555) );
NOR2_X4 U_g24557 ( .A1(g15699), .A2(g23942), .ZN(g24557) );
NOR2_X4 U_g24558 ( .A1(g23917), .A2(g22804), .ZN(g24558) );
NOR2_X4 U_g24566 ( .A1(g23944), .A2(g22842), .ZN(g24566) );
NOR2_X4 U_g24575 ( .A1(g23972), .A2(g22874), .ZN(g24575) );
NOR2_X4 U_g24606 ( .A1(g24183), .A2(g537), .ZN(g24606) );
NOR2_X4 U_g24613 ( .A1(g23592), .A2(g22515), .ZN(g24613) );
NOR2_X4 U_g24622 ( .A1(g23616), .A2(g22546), .ZN(g24622) );
NOR2_X4 U_g24623 ( .A1(g24183), .A2(g529), .ZN(g24623) );
NOR2_X4 U_g24624 ( .A1(g23624), .A2(g22555), .ZN(g24624) );
NOR2_X4 U_g24636 ( .A1(g24183), .A2(g530), .ZN(g24636) );
NOR2_X4 U_g24637 ( .A1(g23665), .A2(g22587), .ZN(g24637) );
NOR2_X4 U_g24638 ( .A1(g23673), .A2(g22595), .ZN(g24638) );
NOR2_X4 U_g24652 ( .A1(g24183), .A2(g531), .ZN(g24652) );
NOR2_X4 U_g24656 ( .A1(g23715), .A2(g22624), .ZN(g24656) );
NOR2_X4 U_g24657 ( .A1(g23723), .A2(g22632), .ZN(g24657) );
NOR2_X4 U_g24663 ( .A1(g24183), .A2(g532), .ZN(g24663) );
NOR2_X4 U_g24675 ( .A1(g23769), .A2(g22660), .ZN(g24675) );
NOR2_X4 U_g24681 ( .A1(g24183), .A2(g533), .ZN(g24681) );
NOR2_X4 U_g24682 ( .A1(g23688), .A2(g24183), .ZN(g24682) );
NOR2_X4 U_g24694 ( .A1(g24183), .A2(g534), .ZN(g24694) );
NOR2_X4 U_g24708 ( .A1(g23854), .A2(g22727), .ZN(g24708) );
NOR2_X4 U_g24711 ( .A1(g24183), .A2(g536), .ZN(g24711) );
NOR2_X4 U_g24717 ( .A1(g23886), .A2(g22754), .ZN(g24717) );
NOR2_X4 U_g24720 ( .A1(g23888), .A2(g22759), .ZN(g24720) );
NOR2_X4 U_g24728 ( .A1(g23907), .A2(g22788), .ZN(g24728) );
NOR2_X4 U_g24731 ( .A1(g23909), .A2(g22793), .ZN(g24731) );
NOR2_X4 U_g24736 ( .A1(g23939), .A2(g22830), .ZN(g24736) );
NOR2_X4 U_g24739 ( .A1(g23941), .A2(g22835), .ZN(g24739) );
NOR2_X4 U_g24742 ( .A1(g23971), .A2(g22869), .ZN(g24742) );
NOR2_X4 U_g24756 ( .A1(g16089), .A2(g24211), .ZN(g24756) );
NOR2_X4 U_g24770 ( .A1(g16119), .A2(g24217), .ZN(g24770) );
NOR2_X4 U_g24782 ( .A1(g16160), .A2(g24221), .ZN(g24782) );
NOR2_X4 U_g24783 ( .A1(g16161), .A2(g24224), .ZN(g24783) );
NOR2_X4 U_g24800 ( .A1(g16211), .A2(g24229), .ZN(g24800) );
NOR2_X4 U_g24819 ( .A1(g16262), .A2(g24236), .ZN(g24819) );
NOR2_X4 U_g24836 ( .A1(g16309), .A2(g24241), .ZN(g24836) );
NOR2_X4 U_g24845 ( .A1(g16350), .A2(g24246), .ZN(g24845) );
NOR2_X4 U_g24847 ( .A1(g16356), .A2(g24247), .ZN(g24847) );
NOR2_X4 U_g24859 ( .A1(g16390), .A2(g24253), .ZN(g24859) );
NOR2_X4 U_g24871 ( .A1(g16422), .A2(g24256), .ZN(g24871) );
NOR2_X4 U_g25027 ( .A1(g24227), .A2(g17001), .ZN(g25027) );
NOR2_X4 U_g25042 ( .A1(g24234), .A2(g17031), .ZN(g25042) );
NOR2_X4 U_g25056 ( .A1(g24242), .A2(g17065), .ZN(g25056) );
NOR2_X4 U_g25067 ( .A1(g24249), .A2(g17100), .ZN(g25067) );
NOR2_X4 U_g25075 ( .A1(g13880), .A2(g23483), .ZN(g25075) );
NOR2_X4 U_g25076 ( .A1(g23409), .A2(g22187), .ZN(g25076) );
NOR2_X4 U_g25077 ( .A1(g23414), .A2(g22196), .ZN(g25077) );
NOR2_X4 U_g25078 ( .A1(g23419), .A2(g22201), .ZN(g25078) );
NOR2_X4 U_g25081 ( .A1(g23423), .A2(g22202), .ZN(g25081) );
NOR2_X4 U_g25082 ( .A1(g23428), .A2(g22207), .ZN(g25082) );
NOR2_X4 U_g25085 ( .A1(g23432), .A2(g22208), .ZN(g25085) );
NOR2_X4 U_g25091 ( .A1(g23434), .A2(g22215), .ZN(g25091) );
NOR2_X4 U_g25099 ( .A1(g23440), .A2(g22224), .ZN(g25099) );
NOR2_X4 U_g25125 ( .A1(g23510), .A2(g22340), .ZN(g25125) );
NOR2_X4 U_g25127 ( .A1(g23525), .A2(g22363), .ZN(g25127) );
NOR2_X4 U_g25129 ( .A1(g23536), .A2(g22383), .ZN(g25129) );
NOR2_X4 U_g25185 ( .A1(g24492), .A2(g10024), .ZN(g25185) );
NOR2_X4 U_g25189 ( .A1(g24502), .A2(g10133), .ZN(g25189) );
NOR2_X4 U_g25191 ( .A1(g24516), .A2(g22777), .ZN(g25191) );
NOR2_X4 U_g25194 ( .A1(g24514), .A2(g10238), .ZN(g25194) );
NOR2_X4 U_g25197 ( .A1(g24528), .A2(g10340), .ZN(g25197) );
NOR2_X4 U_g25199 ( .A1(g24558), .A2(g20127), .ZN(g25199) );
NOR2_X4 U_g25201 ( .A1(g24575), .A2(g18407), .ZN(g25201) );
NOR2_X4 U_g25202 ( .A1(g24566), .A2(g22907), .ZN(g25202) );
NOR2_X4 U_g25204 ( .A1(g24745), .A2(g23547), .ZN(g25204) );
NOR2_X4 U_g25206 ( .A1(g24746), .A2(g23550), .ZN(g25206) );
NOR2_X4 U_g25207 ( .A1(g24747), .A2(g23551), .ZN(g25207) );
NOR2_X4 U_g25208 ( .A1(g24748), .A2(g23552), .ZN(g25208) );
NOR2_X4 U_g25209 ( .A1(g24749), .A2(g23554), .ZN(g25209) );
NOR2_X4 U_g25211 ( .A1(g24750), .A2(g23558), .ZN(g25211) );
NOR2_X4 U_g25212 ( .A1(g24751), .A2(g23559), .ZN(g25212) );
NOR2_X4 U_g25213 ( .A1(g24752), .A2(g23560), .ZN(g25213) );
NOR2_X4 U_g25214 ( .A1(g24754), .A2(g23563), .ZN(g25214) );
NOR2_X4 U_g25215 ( .A1(g24755), .A2(g23564), .ZN(g25215) );
NOR2_X4 U_g25216 ( .A1(g24757), .A2(g23565), .ZN(g25216) );
NOR2_X4 U_g25217 ( .A1(g24758), .A2(g23567), .ZN(g25217) );
NOR2_X4 U_g25218 ( .A1(g24760), .A2(g23571), .ZN(g25218) );
NOR2_X4 U_g25219 ( .A1(g24761), .A2(g23572), .ZN(g25219) );
NOR2_X4 U_g25220 ( .A1(g24762), .A2(g23573), .ZN(g25220) );
NOR2_X4 U_g25221 ( .A1(g24767), .A2(g23577), .ZN(g25221) );
NOR2_X4 U_g25222 ( .A1(g24768), .A2(g23578), .ZN(g25222) );
NOR2_X4 U_g25223 ( .A1(g24769), .A2(g23579), .ZN(g25223) );
NOR2_X4 U_g25224 ( .A1(g24772), .A2(g23582), .ZN(g25224) );
NOR2_X4 U_g25225 ( .A1(g24773), .A2(g23583), .ZN(g25225) );
NOR2_X4 U_g25226 ( .A1(g24774), .A2(g23584), .ZN(g25226) );
NOR2_X4 U_g25227 ( .A1(g24775), .A2(g23586), .ZN(g25227) );
NOR2_X4 U_g25228 ( .A1(g24776), .A2(g23590), .ZN(g25228) );
NOR2_X4 U_g25229 ( .A1(g24777), .A2(g23591), .ZN(g25229) );
NOR2_X4 U_g25230 ( .A1(g24779), .A2(g23598), .ZN(g25230) );
NOR2_X4 U_g25231 ( .A1(g24780), .A2(g23599), .ZN(g25231) );
NOR2_X4 U_g25232 ( .A1(g24781), .A2(g23600), .ZN(g25232) );
NOR2_X4 U_g25233 ( .A1(g24788), .A2(g23604), .ZN(g25233) );
NOR2_X4 U_g25234 ( .A1(g24789), .A2(g23605), .ZN(g25234) );
NOR2_X4 U_g25235 ( .A1(g24790), .A2(g23606), .ZN(g25235) );
NOR2_X4 U_g25236 ( .A1(g24792), .A2(g23609), .ZN(g25236) );
NOR2_X4 U_g25237 ( .A1(g24793), .A2(g23610), .ZN(g25237) );
NOR2_X4 U_g25238 ( .A1(g24794), .A2(g23611), .ZN(g25238) );
NOR2_X4 U_g25239 ( .A1(g24796), .A2(g23615), .ZN(g25239) );
NOR2_X4 U_g25240 ( .A1(g24798), .A2(g23622), .ZN(g25240) );
NOR2_X4 U_g25241 ( .A1(g24799), .A2(g23623), .ZN(g25241) );
NOR2_X4 U_g25242 ( .A1(g24802), .A2(g23630), .ZN(g25242) );
NOR2_X4 U_g25243 ( .A1(g24803), .A2(g23631), .ZN(g25243) );
NOR2_X4 U_g25244 ( .A1(g24804), .A2(g23632), .ZN(g25244) );
NOR2_X4 U_g25245 ( .A1(g24809), .A2(g23636), .ZN(g25245) );
NOR2_X4 U_g25246 ( .A1(g24810), .A2(g23637), .ZN(g25246) );
NOR2_X4 U_g25247 ( .A1(g24811), .A2(g23638), .ZN(g25247) );
NOR2_X4 U_g25248 ( .A1(g24818), .A2(g23664), .ZN(g25248) );
NOR2_X4 U_g25249 ( .A1(g24821), .A2(g23671), .ZN(g25249) );
NOR2_X4 U_g25250 ( .A1(g24822), .A2(g23672), .ZN(g25250) );
NOR2_X4 U_g25251 ( .A1(g24824), .A2(g23679), .ZN(g25251) );
NOR2_X4 U_g25252 ( .A1(g24825), .A2(g23680), .ZN(g25252) );
NOR2_X4 U_g25253 ( .A1(g24826), .A2(g23681), .ZN(g25253) );
NOR2_X4 U_g25254 ( .A1(g24831), .A2(g23687), .ZN(g25254) );
NOR2_X4 U_g25255 ( .A1(g24838), .A2(g23714), .ZN(g25255) );
NOR2_X4 U_g25256 ( .A1(g24840), .A2(g23721), .ZN(g25256) );
NOR2_X4 U_g25257 ( .A1(g24841), .A2(g23722), .ZN(g25257) );
NOR2_X4 U_g25258 ( .A1(g24846), .A2(g23741), .ZN(g25258) );
NOR2_X4 U_g25259 ( .A1(g24853), .A2(g23768), .ZN(g25259) );
NOR2_X4 U_g25260 ( .A1(g24858), .A2(g17737), .ZN(g25260) );
NOR2_X4 U_g25261 ( .A1(g24861), .A2(g23796), .ZN(g25261) );
NOR2_X4 U_g25262 ( .A1(g24869), .A2(g17824), .ZN(g25262) );
NOR2_X4 U_g25263 ( .A1(g24874), .A2(g17838), .ZN(g25263) );
NOR2_X4 U_g25264 ( .A1(g24876), .A2(g23849), .ZN(g25264) );
NOR2_X4 U_g25265 ( .A1(g24878), .A2(g23852), .ZN(g25265) );
NOR2_X4 U_g25266 ( .A1(g24881), .A2(g17912), .ZN(g25266) );
NOR2_X4 U_g25267 ( .A1(g24884), .A2(g17936), .ZN(g25267) );
NOR2_X4 U_g25268 ( .A1(g24888), .A2(g17950), .ZN(g25268) );
NOR2_X4 U_g25270 ( .A1(g24898), .A2(g18023), .ZN(g25270) );
NOR2_X4 U_g25271 ( .A1(g24901), .A2(g18047), .ZN(g25271) );
NOR2_X4 U_g25272 ( .A1(g24905), .A2(g18061), .ZN(g25272) );
NOR2_X4 U_g25273 ( .A1(g24907), .A2(g23904), .ZN(g25273) );
NOR2_X4 U_g25279 ( .A1(g24921), .A2(g18140), .ZN(g25279) );
NOR2_X4 U_g25280 ( .A1(g24924), .A2(g18164), .ZN(g25280) );
NOR2_X4 U_g25288 ( .A1(g24938), .A2(g18256), .ZN(g25288) );
NOR2_X4 U_g25311 ( .A1(g24964), .A2(g24029), .ZN(g25311) );
NOR2_X4 U_g25343 ( .A1(g24975), .A2(g5623), .ZN(g25343) );
NOR2_X4 U_g25357 ( .A1(g24986), .A2(g5651), .ZN(g25357) );
NOR2_X4 U_g25372 ( .A1(g24997), .A2(g5689), .ZN(g25372) );
NOR2_X4 U_g25389 ( .A1(g25005), .A2(g5741), .ZN(g25389) );
NOR2_X4 U_g25418 ( .A1(g24482), .A2(g22319), .ZN(g25418) );
NOR2_X4 U_g25426 ( .A1(g24183), .A2(g24616), .ZN(g25426) );
NOR2_X4 U_g25429 ( .A1(g24482), .A2(g22319), .ZN(g25429) );
NOR2_X4 U_g25450 ( .A1(g16018), .A2(g25086), .ZN(g25450) );
NOR2_X4 U_g25451 ( .A1(g16048), .A2(g25102), .ZN(g25451) );
NOR2_X4 U_g25452 ( .A1(g16101), .A2(g25117), .ZN(g25452) );
NOR2_X4 U_g25523 ( .A1(g20842), .A2(g24429), .ZN(g25523) );
NOR2_X4 U_g25539 ( .A1(g25088), .A2(g6157), .ZN(g25539) );
NOR2_X4 U_g25569 ( .A1(g24708), .A2(g24490), .ZN(g25569) );
NOR2_X4 U_g25589 ( .A1(g20850), .A2(g24433), .ZN(g25589) );
NOR2_X4 U_g25605 ( .A1(g25096), .A2(g6184), .ZN(g25605) );
NOR2_X4 U_g25631 ( .A1(g24717), .A2(g24497), .ZN(g25631) );
NOR2_X4 U_g25648 ( .A1(g24720), .A2(g24500), .ZN(g25648) );
NOR2_X4 U_g25668 ( .A1(g20858), .A2(g24437), .ZN(g25668) );
NOR2_X4 U_g25684 ( .A1(g25106), .A2(g6216), .ZN(g25684) );
NOR2_X4 U_g25699 ( .A1(g24613), .A2(g24506), .ZN(g25699) );
NOR2_X4 U_g25708 ( .A1(g24728), .A2(g24509), .ZN(g25708) );
NOR2_X4 U_g25725 ( .A1(g24731), .A2(g24512), .ZN(g25725) );
NOR2_X4 U_g25745 ( .A1(g20866), .A2(g24440), .ZN(g25745) );
NOR2_X4 U_g25761 ( .A1(g25112), .A2(g6305), .ZN(g25761) );
NOR2_X4 U_g25764 ( .A1(g25076), .A2(g21615), .ZN(g25764) );
NOR2_X4 U_g25772 ( .A1(g24624), .A2(g24520), .ZN(g25772) );
NOR2_X4 U_g25781 ( .A1(g24736), .A2(g24523), .ZN(g25781) );
NOR2_X4 U_g25798 ( .A1(g24739), .A2(g24526), .ZN(g25798) );
NOR2_X4 U_g25818 ( .A1(g25077), .A2(g21643), .ZN(g25818) );
NOR2_X4 U_g25826 ( .A1(g24638), .A2(g24533), .ZN(g25826) );
NOR2_X4 U_g25835 ( .A1(g24742), .A2(g24536), .ZN(g25835) );
NOR3_X4 U_g25852 ( .A1(g4456), .A2(g14831), .A3(g25078), .ZN(g25852) );
NOR2_X4 U_g25853 ( .A1(g25081), .A2(g21674), .ZN(g25853) );
NOR2_X4 U_g25861 ( .A1(g24657), .A2(g24546), .ZN(g25861) );
NOR4_X4 U_g25870 ( .A1(g4456), .A2(g25078), .A3(g18429), .A4(g16075), .ZN(g25870) );
NOR3_X4 U_g25873 ( .A1(g4632), .A2(g14904), .A3(g25082), .ZN(g25873) );
NOR2_X4 U_g25874 ( .A1(g25085), .A2(g21703), .ZN(g25874) );
NOR4_X4 U_g25882 ( .A1(g4632), .A2(g25082), .A3(g18502), .A4(g16113), .ZN(g25882) );
NOR3_X4 U_g25885 ( .A1(g4809), .A2(g14985), .A3(g25091), .ZN(g25885) );
NOR4_X4 U_g25887 ( .A1(g4809), .A2(g25091), .A3(g18566), .A4(g16164), .ZN(g25887) );
NOR3_X4 U_g25890 ( .A1(g4985), .A2(g15074), .A3(g25099), .ZN(g25890) );
NOR4_X4 U_g25892 ( .A1(g4985), .A2(g25099), .A3(g18616), .A4(g16223), .ZN(g25892) );
NOR2_X4 U_g25932 ( .A1(g25125), .A2(g17001), .ZN(g25932) );
NOR2_X4 U_g25935 ( .A1(g25127), .A2(g17031), .ZN(g25935) );
NOR2_X4 U_g25938 ( .A1(g25129), .A2(g17065), .ZN(g25938) );
NOR2_X4 U_g25940 ( .A1(g24428), .A2(g17100), .ZN(g25940) );
NOR2_X4 U_g25941 ( .A1(g24529), .A2(g24540), .ZN(g25941) );
NOR2_X4 U_g25943 ( .A1(g24541), .A2(g24550), .ZN(g25943) );
NOR2_X4 U_g25944 ( .A1(g24542), .A2(g24552), .ZN(g25944) );
NOR2_X4 U_g25946 ( .A1(g24553), .A2(g24561), .ZN(g25946) );
NOR2_X4 U_g25947 ( .A1(g24554), .A2(g24563), .ZN(g25947) );
NOR2_X4 U_g25948 ( .A1(g24564), .A2(g24571), .ZN(g25948) );
NOR2_X4 U_g25949 ( .A1(g24565), .A2(g24573), .ZN(g25949) );
NOR2_X4 U_g25950 ( .A1(g24574), .A2(g24580), .ZN(g25950) );
NOR2_X4 U_g25962 ( .A1(g24591), .A2(g23496), .ZN(g25962) );
NOR2_X4 U_g25967 ( .A1(g24596), .A2(g23512), .ZN(g25967) );
NOR2_X4 U_g25974 ( .A1(g24604), .A2(g23527), .ZN(g25974) );
NOR2_X4 U_g25979 ( .A1(g24611), .A2(g23538), .ZN(g25979) );
NOR2_X4 U_g26025 ( .A1(g25392), .A2(g17193), .ZN(g26025) );
NOR2_X4 U_g26031 ( .A1(g25273), .A2(g22777), .ZN(g26031) );
NOR2_X4 U_g26037 ( .A1(g25311), .A2(g18407), .ZN(g26037) );
NOR2_X4 U_g26041 ( .A1(g25475), .A2(g24855), .ZN(g26041) );
NOR2_X4 U_g26042 ( .A1(g25505), .A2(g24867), .ZN(g26042) );
NOR2_X4 U_g26043 ( .A1(g25506), .A2(g24870), .ZN(g26043) );
NOR2_X4 U_g26044 ( .A1(g25552), .A2(g24882), .ZN(g26044) );
NOR2_X4 U_g26045 ( .A1(g25553), .A2(g24885), .ZN(g26045) );
NOR2_X4 U_g26046 ( .A1(g25618), .A2(g24899), .ZN(g26046) );
NOR2_X4 U_g26047 ( .A1(g25619), .A2(g24902), .ZN(g26047) );
NOR2_X4 U_g26048 ( .A1(g25628), .A2(g24906), .ZN(g26048) );
NOR2_X4 U_g26049 ( .A1(g25629), .A2(g24908), .ZN(g26049) );
NOR2_X4 U_g26050 ( .A1(g25697), .A2(g24922), .ZN(g26050) );
NOR2_X4 U_g26055 ( .A1(g25881), .A2(g24974), .ZN(g26055) );
NOR2_X4 U_g26081 ( .A1(g25470), .A2(g25482), .ZN(g26081) );
NOR2_X4 U_g26083 ( .A1(g25426), .A2(g22319), .ZN(g26083) );
NOR2_X4 U_g26084 ( .A1(g25487), .A2(g25513), .ZN(g26084) );
NOR3_X4 U_g26087 ( .A1(g6068), .A2(g24183), .A3(g25319), .ZN(g26087) );
NOR2_X4 U_g26090 ( .A1(g25518), .A2(g25560), .ZN(g26090) );
NOR3_X4 U_g26096 ( .A1(g6068), .A2(g24183), .A3(g25394), .ZN(g26096) );
NOR3_X4 U_g26099 ( .A1(g6068), .A2(g24183), .A3(g25313), .ZN(g26099) );
NOR2_X4 U_g26103 ( .A1(g25565), .A2(g25626), .ZN(g26103) );
NOR3_X4 U_g26107 ( .A1(g6068), .A2(g24183), .A3(g25383), .ZN(g26107) );
NOR3_X4 U_g26110 ( .A1(g6068), .A2(g24183), .A3(g25305), .ZN(g26110) );
NOR2_X4 U_g26113 ( .A1(g25426), .A2(g22319), .ZN(g26113) );
NOR3_X4 U_g26126 ( .A1(g6068), .A2(g24183), .A3(g25368), .ZN(g26126) );
NOR3_X4 U_g26137 ( .A1(g6068), .A2(g24183), .A3(g25355), .ZN(g26137) );
NOR2_X4 U_g26140 ( .A1(g24183), .A2(g25430), .ZN(g26140) );
NOR3_X4 U_g26145 ( .A1(g6068), .A2(g24183), .A3(g25347), .ZN(g26145) );
NOR3_X4 U_g26151 ( .A1(g6068), .A2(g24183), .A3(g25335), .ZN(g26151) );
NOR3_X4 U_g26154 ( .A1(g6068), .A2(g24183), .A3(g25329), .ZN(g26154) );
NOR2_X4 U_g26160 ( .A1(g25951), .A2(g16162), .ZN(g26160) );
NOR2_X4 U_g26168 ( .A1(g25953), .A2(g16212), .ZN(g26168) );
NOR2_X4 U_g26183 ( .A1(g25957), .A2(g13270), .ZN(g26183) );
NOR2_X4 U_g26199 ( .A1(g25961), .A2(g13291), .ZN(g26199) );
NOR2_X4 U_g26217 ( .A1(g25963), .A2(g13320), .ZN(g26217) );
NOR2_X4 U_g26240 ( .A1(g25968), .A2(g13340), .ZN(g26240) );
NOR2_X4 U_g26265 ( .A1(g25972), .A2(g13360), .ZN(g26265) );
NOR2_X4 U_g26272 ( .A1(g25973), .A2(g16423), .ZN(g26272) );
NOR2_X4 U_g26283 ( .A1(g25954), .A2(g24486), .ZN(g26283) );
NOR2_X4 U_g26295 ( .A1(g25977), .A2(g13385), .ZN(g26295) );
NOR2_X4 U_g26304 ( .A1(g25978), .A2(g16451), .ZN(g26304) );
NOR2_X4 U_g26327 ( .A1(g25958), .A2(g24493), .ZN(g26327) );
NOR2_X4 U_g26336 ( .A1(g25981), .A2(g13481), .ZN(g26336) );
NOR2_X4 U_g26374 ( .A1(g25964), .A2(g24503), .ZN(g26374) );
NOR2_X4 U_g26417 ( .A1(g25969), .A2(g24515), .ZN(g26417) );
NOR2_X4 U_g26529 ( .A1(g25962), .A2(g17001), .ZN(g26529) );
NOR2_X4 U_g26530 ( .A1(g25967), .A2(g17031), .ZN(g26530) );
NOR2_X4 U_g26531 ( .A1(g25974), .A2(g17065), .ZN(g26531) );
NOR2_X4 U_g26532 ( .A1(g25979), .A2(g17100), .ZN(g26532) );
NOR2_X4 U_g26534 ( .A1(g25321), .A2(g8869), .ZN(g26534) );
NOR2_X4 U_g26541 ( .A1(g13755), .A2(g25269), .ZN(g26541) );
NOR2_X4 U_g26545 ( .A1(g13790), .A2(g25277), .ZN(g26545) );
NOR2_X4 U_g26547 ( .A1(g13796), .A2(g25278), .ZN(g26547) );
NOR2_X4 U_g26553 ( .A1(g13816), .A2(g25282), .ZN(g26553) );
NOR2_X4 U_g26557 ( .A1(g13818), .A2(g25286), .ZN(g26557) );
NOR2_X4 U_g26559 ( .A1(g13824), .A2(g25287), .ZN(g26559) );
NOR2_X4 U_g26560 ( .A1(g25281), .A2(g24559), .ZN(g26560) );
NOR2_X4 U_g26569 ( .A1(g13837), .A2(g25290), .ZN(g26569) );
NOR2_X4 U_g26573 ( .A1(g13839), .A2(g25294), .ZN(g26573) );
NOR2_X4 U_g26575 ( .A1(g13845), .A2(g25295), .ZN(g26575) );
NOR2_X4 U_g26583 ( .A1(g25289), .A2(g24569), .ZN(g26583) );
NOR2_X4 U_g26592 ( .A1(g13851), .A2(g25300), .ZN(g26592) );
NOR2_X4 U_g26596 ( .A1(g13853), .A2(g25304), .ZN(g26596) );
NOR2_X4 U_g26607 ( .A1(g25299), .A2(g24578), .ZN(g26607) );
NOR2_X4 U_g26616 ( .A1(g13860), .A2(g25310), .ZN(g26616) );
NOR2_X4 U_g26630 ( .A1(g25309), .A2(g24585), .ZN(g26630) );
NOR2_X4 U_g26655 ( .A1(g25328), .A2(g17084), .ZN(g26655) );
NOR2_X4 U_g26659 ( .A1(g25334), .A2(g17116), .ZN(g26659) );
NOR2_X4 U_g26660 ( .A1(g25208), .A2(g10024), .ZN(g26660) );
NOR2_X4 U_g26661 ( .A1(g25337), .A2(g17122), .ZN(g26661) );
NOR2_X4 U_g26664 ( .A1(g25346), .A2(g17138), .ZN(g26664) );
NOR2_X4 U_g26665 ( .A1(g25348), .A2(g17143), .ZN(g26665) );
NOR2_X4 U_g26666 ( .A1(g25216), .A2(g10133), .ZN(g26666) );
NOR2_X4 U_g26667 ( .A1(g25351), .A2(g17149), .ZN(g26667) );
NOR2_X4 U_g26669 ( .A1(g25360), .A2(g17161), .ZN(g26669) );
NOR2_X4 U_g26670 ( .A1(g25362), .A2(g17166), .ZN(g26670) );
NOR2_X4 U_g26671 ( .A1(g25226), .A2(g10238), .ZN(g26671) );
NOR2_X4 U_g26672 ( .A1(g25365), .A2(g17172), .ZN(g26672) );
NOR2_X4 U_g26675 ( .A1(g25375), .A2(g17176), .ZN(g26675) );
NOR2_X4 U_g26676 ( .A1(g25377), .A2(g17181), .ZN(g26676) );
NOR2_X4 U_g26677 ( .A1(g25238), .A2(g10340), .ZN(g26677) );
NOR2_X4 U_g26776 ( .A1(g26042), .A2(g10024), .ZN(g26776) );
NOR2_X4 U_g26781 ( .A1(g26044), .A2(g10133), .ZN(g26781) );
NOR2_X4 U_g26786 ( .A1(g26049), .A2(g22777), .ZN(g26786) );
NOR2_X4 U_g26789 ( .A1(g26046), .A2(g10238), .ZN(g26789) );
NOR2_X4 U_g26795 ( .A1(g26050), .A2(g10340), .ZN(g26795) );
NOR2_X4 U_g26798 ( .A1(g26055), .A2(g18407), .ZN(g26798) );
NOR2_X4 U_g26799 ( .A1(g26158), .A2(g25453), .ZN(g26799) );
NOR2_X4 U_g26800 ( .A1(g26163), .A2(g25457), .ZN(g26800) );
NOR2_X4 U_g26801 ( .A1(g26171), .A2(g25461), .ZN(g26801) );
NOR2_X4 U_g26802 ( .A1(g26188), .A2(g25466), .ZN(g26802) );
NOR2_X4 U_g26803 ( .A1(g15105), .A2(g26213), .ZN(g26803) );
NOR2_X4 U_g26804 ( .A1(g15172), .A2(g26235), .ZN(g26804) );
NOR2_X4 U_g26805 ( .A1(g15173), .A2(g26236), .ZN(g26805) );
NOR2_X4 U_g26806 ( .A1(g15197), .A2(g26244), .ZN(g26806) );
NOR2_X4 U_g26807 ( .A1(g15245), .A2(g26261), .ZN(g26807) );
NOR2_X4 U_g26808 ( .A1(g15246), .A2(g26262), .ZN(g26808) );
NOR2_X4 U_g26809 ( .A1(g15258), .A2(g26270), .ZN(g26809) );
NOR2_X4 U_g26810 ( .A1(g15259), .A2(g26271), .ZN(g26810) );
NOR2_X4 U_g26811 ( .A1(g15283), .A2(g26279), .ZN(g26811) );
NOR2_X4 U_g26812 ( .A1(g15321), .A2(g26291), .ZN(g26812) );
NOR2_X4 U_g26813 ( .A1(g15337), .A2(g26302), .ZN(g26813) );
NOR2_X4 U_g26814 ( .A1(g15338), .A2(g26303), .ZN(g26814) );
NOR2_X4 U_g26815 ( .A1(g15350), .A2(g26311), .ZN(g26815) );
NOR2_X4 U_g26816 ( .A1(g15351), .A2(g26312), .ZN(g26816) );
NOR2_X4 U_g26817 ( .A1(g15375), .A2(g26317), .ZN(g26817) );
NOR2_X4 U_g26818 ( .A1(g15407), .A2(g26335), .ZN(g26818) );
NOR2_X4 U_g26820 ( .A1(g15423), .A2(g26346), .ZN(g26820) );
NOR2_X4 U_g26821 ( .A1(g15424), .A2(g26347), .ZN(g26821) );
NOR2_X4 U_g26822 ( .A1(g15436), .A2(g26352), .ZN(g26822) );
NOR2_X4 U_g26823 ( .A1(g15437), .A2(g26353), .ZN(g26823) );
NOR2_X4 U_g26824 ( .A1(g15491), .A2(g26382), .ZN(g26824) );
NOR2_X4 U_g26825 ( .A1(g15507), .A2(g26390), .ZN(g26825) );
NOR2_X4 U_g26826 ( .A1(g15508), .A2(g26391), .ZN(g26826) );
NOR2_X4 U_g26827 ( .A1(g15577), .A2(g26425), .ZN(g26827) );
NOR2_X4 U_g26869 ( .A1(g26458), .A2(g5642), .ZN(g26869) );
NOR2_X4 U_g26873 ( .A1(g25483), .A2(g26260), .ZN(g26873) );
NOR2_X4 U_g26877 ( .A1(g26140), .A2(g22319), .ZN(g26877) );
NOR2_X4 U_g26878 ( .A1(g26482), .A2(g5680), .ZN(g26878) );
NOR2_X4 U_g26882 ( .A1(g25514), .A2(g26301), .ZN(g26882) );
NOR2_X4 U_g26885 ( .A1(g26140), .A2(g22319), .ZN(g26885) );
NOR2_X4 U_g26887 ( .A1(g26498), .A2(g5732), .ZN(g26887) );
NOR2_X4 U_g26891 ( .A1(g25561), .A2(g26345), .ZN(g26891) );
NOR2_X4 U_g26897 ( .A1(g26513), .A2(g5790), .ZN(g26897) );
NOR2_X4 U_g26901 ( .A1(g25627), .A2(g26389), .ZN(g26901) );
NOR2_X4 U_g26905 ( .A1(g26096), .A2(g22319), .ZN(g26905) );
NOR2_X4 U_g26914 ( .A1(g26107), .A2(g22319), .ZN(g26914) );
NOR2_X4 U_g26988 ( .A1(g24893), .A2(g26023), .ZN(g26988) );
NOR2_X4 U_g26989 ( .A1(g26663), .A2(g21913), .ZN(g26989) );
NOR2_X4 U_g27011 ( .A1(g24916), .A2(g26026), .ZN(g27011) );
NOR2_X4 U_g27012 ( .A1(g26668), .A2(g21931), .ZN(g27012) );
NOR2_X4 U_g27037 ( .A1(g24933), .A2(g26028), .ZN(g27037) );
NOR2_X4 U_g27038 ( .A1(g26674), .A2(g20640), .ZN(g27038) );
NOR2_X4 U_g27051 ( .A1(g4456), .A2(g26081), .ZN(g27051) );
NOR2_X4 U_g27065 ( .A1(g24945), .A2(g26029), .ZN(g27065) );
NOR2_X4 U_g27066 ( .A1(g26024), .A2(g20665), .ZN(g27066) );
NOR2_X4 U_g27078 ( .A1(g4632), .A2(g26084), .ZN(g27078) );
NOR2_X4 U_g27094 ( .A1(g4809), .A2(g26090), .ZN(g27094) );
NOR2_X4 U_g27106 ( .A1(g4985), .A2(g26103), .ZN(g27106) );
NOR2_X4 U_g27120 ( .A1(g26560), .A2(g17001), .ZN(g27120) );
NOR2_X4 U_g27123 ( .A1(g26583), .A2(g17031), .ZN(g27123) );
NOR2_X4 U_g27129 ( .A1(g26607), .A2(g17065), .ZN(g27129) );
NOR2_X4 U_g27131 ( .A1(g26630), .A2(g17100), .ZN(g27131) );
NOR2_X4 U_g27144 ( .A1(g23451), .A2(g26052), .ZN(g27144) );
NOR2_X4 U_g27147 ( .A1(g23458), .A2(g26054), .ZN(g27147) );
NOR2_X4 U_g27149 ( .A1(g23462), .A2(g26060), .ZN(g27149) );
NOR2_X4 U_g27152 ( .A1(g23467), .A2(g26062), .ZN(g27152) );
NOR2_X4 U_g27157 ( .A1(g23471), .A2(g26067), .ZN(g27157) );
NOR2_X4 U_g27160 ( .A1(g23476), .A2(g26069), .ZN(g27160) );
NOR2_X4 U_g27165 ( .A1(g23484), .A2(g26074), .ZN(g27165) );
NOR2_X4 U_g27174 ( .A1(g23494), .A2(g26080), .ZN(g27174) );
NOR2_X4 U_g27175 ( .A1(g26075), .A2(g25342), .ZN(g27175) );
NOR2_X4 U_g27179 ( .A1(g26082), .A2(g25356), .ZN(g27179) );
NOR2_X4 U_g27184 ( .A1(g26085), .A2(g25371), .ZN(g27184) );
NOR2_X4 U_g27188 ( .A1(g26091), .A2(g25388), .ZN(g27188) );
NOR2_X4 U_g27243 ( .A1(g26802), .A2(g10340), .ZN(g27243) );
NOR2_X4 U_g27250 ( .A1(g26955), .A2(g26166), .ZN(g27250) );
NOR2_X4 U_g27251 ( .A1(g26958), .A2(g26186), .ZN(g27251) );
NOR2_X4 U_g27252 ( .A1(g26963), .A2(g26207), .ZN(g27252) );
NOR2_X4 U_g27253 ( .A1(g26965), .A2(g26212), .ZN(g27253) );
NOR2_X4 U_g27254 ( .A1(g26968), .A2(g26231), .ZN(g27254) );
NOR2_X4 U_g27255 ( .A1(g26969), .A2(g26233), .ZN(g27255) );
NOR2_X4 U_g27256 ( .A1(g26970), .A2(g26234), .ZN(g27256) );
NOR2_X4 U_g27257 ( .A1(g26971), .A2(g26243), .ZN(g27257) );
NOR2_X4 U_g27258 ( .A1(g26977), .A2(g26257), .ZN(g27258) );
NOR2_X4 U_g27259 ( .A1(g26978), .A2(g26258), .ZN(g27259) );
NOR2_X4 U_g27260 ( .A1(g26979), .A2(g26259), .ZN(g27260) );
NOR2_X4 U_g27261 ( .A1(g26980), .A2(g26263), .ZN(g27261) );
NOR2_X4 U_g27262 ( .A1(g26981), .A2(g26268), .ZN(g27262) );
NOR2_X4 U_g27263 ( .A1(g26982), .A2(g26269), .ZN(g27263) );
NOR2_X4 U_g27264 ( .A1(g26984), .A2(g26278), .ZN(g27264) );
NOR2_X4 U_g27265 ( .A1(g26993), .A2(g26288), .ZN(g27265) );
NOR2_X4 U_g27266 ( .A1(g26994), .A2(g26289), .ZN(g27266) );
NOR2_X4 U_g27267 ( .A1(g26995), .A2(g26290), .ZN(g27267) );
NOR2_X4 U_g27268 ( .A1(g26996), .A2(g26292), .ZN(g27268) );
NOR2_X4 U_g27269 ( .A1(g26997), .A2(g26293), .ZN(g27269) );
NOR2_X4 U_g27270 ( .A1(g26998), .A2(g26298), .ZN(g27270) );
NOR2_X4 U_g27271 ( .A1(g26999), .A2(g26299), .ZN(g27271) );
NOR2_X4 U_g27272 ( .A1(g27000), .A2(g26300), .ZN(g27272) );
NOR2_X4 U_g27273 ( .A1(g27001), .A2(g26307), .ZN(g27273) );
NOR2_X4 U_g27274 ( .A1(g27002), .A2(g26309), .ZN(g27274) );
NOR2_X4 U_g27275 ( .A1(g27003), .A2(g26310), .ZN(g27275) );
NOR2_X4 U_g27276 ( .A1(g27004), .A2(g26316), .ZN(g27276) );
NOR2_X4 U_g27277 ( .A1(g27005), .A2(g26318), .ZN(g27277) );
NOR2_X4 U_g27278 ( .A1(g27006), .A2(g26319), .ZN(g27278) );
NOR2_X4 U_g27279 ( .A1(g27007), .A2(g26324), .ZN(g27279) );
NOR2_X4 U_g27280 ( .A1(g27008), .A2(g26325), .ZN(g27280) );
NOR2_X4 U_g27281 ( .A1(g27009), .A2(g26326), .ZN(g27281) );
NOR2_X4 U_g27282 ( .A1(g27016), .A2(g26332), .ZN(g27282) );
NOR2_X4 U_g27283 ( .A1(g27017), .A2(g26333), .ZN(g27283) );
NOR2_X4 U_g27284 ( .A1(g27018), .A2(g26334), .ZN(g27284) );
NOR2_X4 U_g27285 ( .A1(g27019), .A2(g26339), .ZN(g27285) );
NOR2_X4 U_g27286 ( .A1(g27020), .A2(g26340), .ZN(g27286) );
NOR2_X4 U_g27287 ( .A1(g27021), .A2(g26342), .ZN(g27287) );
NOR2_X4 U_g27288 ( .A1(g27022), .A2(g26343), .ZN(g27288) );
NOR2_X4 U_g27289 ( .A1(g27023), .A2(g26344), .ZN(g27289) );
NOR2_X4 U_g27290 ( .A1(g27024), .A2(g26348), .ZN(g27290) );
NOR2_X4 U_g27291 ( .A1(g27025), .A2(g26350), .ZN(g27291) );
NOR2_X4 U_g27292 ( .A1(g27026), .A2(g26351), .ZN(g27292) );
NOR2_X4 U_g27293 ( .A1(g27027), .A2(g26357), .ZN(g27293) );
NOR2_X4 U_g27294 ( .A1(g27028), .A2(g26361), .ZN(g27294) );
NOR2_X4 U_g27295 ( .A1(g27029), .A2(g26362), .ZN(g27295) );
NOR2_X4 U_g27296 ( .A1(g27030), .A2(g26363), .ZN(g27296) );
NOR2_X4 U_g27297 ( .A1(g27031), .A2(g26365), .ZN(g27297) );
NOR2_X4 U_g27298 ( .A1(g27032), .A2(g26366), .ZN(g27298) );
NOR2_X4 U_g27299 ( .A1(g27033), .A2(g26371), .ZN(g27299) );
NOR2_X4 U_g27300 ( .A1(g27034), .A2(g26372), .ZN(g27300) );
NOR2_X4 U_g27301 ( .A1(g27035), .A2(g26373), .ZN(g27301) );
NOR2_X4 U_g27302 ( .A1(g27042), .A2(g26379), .ZN(g27302) );
NOR2_X4 U_g27303 ( .A1(g27043), .A2(g26380), .ZN(g27303) );
NOR2_X4 U_g27304 ( .A1(g27044), .A2(g26381), .ZN(g27304) );
NOR2_X4 U_g27305 ( .A1(g27045), .A2(g26383), .ZN(g27305) );
NOR2_X4 U_g27306 ( .A1(g27046), .A2(g26384), .ZN(g27306) );
NOR2_X4 U_g27307 ( .A1(g27047), .A2(g26386), .ZN(g27307) );
NOR2_X4 U_g27308 ( .A1(g27048), .A2(g26387), .ZN(g27308) );
NOR2_X4 U_g27309 ( .A1(g27049), .A2(g26388), .ZN(g27309) );
NOR2_X4 U_g27310 ( .A1(g27050), .A2(g26392), .ZN(g27310) );
NOR2_X4 U_g27311 ( .A1(g27053), .A2(g26396), .ZN(g27311) );
NOR2_X4 U_g27312 ( .A1(g27054), .A2(g26397), .ZN(g27312) );
NOR2_X4 U_g27313 ( .A1(g27055), .A2(g26400), .ZN(g27313) );
NOR2_X4 U_g27314 ( .A1(g27056), .A2(g26404), .ZN(g27314) );
NOR2_X4 U_g27315 ( .A1(g27057), .A2(g26405), .ZN(g27315) );
NOR2_X4 U_g27316 ( .A1(g27058), .A2(g26406), .ZN(g27316) );
NOR2_X4 U_g27317 ( .A1(g27059), .A2(g26408), .ZN(g27317) );
NOR2_X4 U_g27318 ( .A1(g27060), .A2(g26409), .ZN(g27318) );
NOR2_X4 U_g27319 ( .A1(g27061), .A2(g26414), .ZN(g27319) );
NOR2_X4 U_g27320 ( .A1(g27062), .A2(g26415), .ZN(g27320) );
NOR2_X4 U_g27321 ( .A1(g27063), .A2(g26416), .ZN(g27321) );
NOR2_X4 U_g27322 ( .A1(g27070), .A2(g26422), .ZN(g27322) );
NOR2_X4 U_g27323 ( .A1(g27071), .A2(g26423), .ZN(g27323) );
NOR2_X4 U_g27324 ( .A1(g27072), .A2(g26424), .ZN(g27324) );
NOR2_X4 U_g27325 ( .A1(g27073), .A2(g26426), .ZN(g27325) );
NOR2_X4 U_g27326 ( .A1(g27074), .A2(g26427), .ZN(g27326) );
NOR2_X4 U_g27327 ( .A1(g27077), .A2(g26432), .ZN(g27327) );
NOR2_X4 U_g27328 ( .A1(g27080), .A2(g26437), .ZN(g27328) );
NOR2_X4 U_g27329 ( .A1(g27081), .A2(g26438), .ZN(g27329) );
NOR2_X4 U_g27330 ( .A1(g27082), .A2(g26441), .ZN(g27330) );
NOR2_X4 U_g27331 ( .A1(g27083), .A2(g26445), .ZN(g27331) );
NOR2_X4 U_g27332 ( .A1(g27084), .A2(g26446), .ZN(g27332) );
NOR2_X4 U_g27333 ( .A1(g27085), .A2(g26447), .ZN(g27333) );
NOR2_X4 U_g27334 ( .A1(g27086), .A2(g26449), .ZN(g27334) );
NOR2_X4 U_g27335 ( .A1(g27087), .A2(g26450), .ZN(g27335) );
NOR2_X4 U_g27336 ( .A1(g27088), .A2(g26455), .ZN(g27336) );
NOR2_X4 U_g27337 ( .A1(g27089), .A2(g26456), .ZN(g27337) );
NOR2_X4 U_g27338 ( .A1(g27090), .A2(g26457), .ZN(g27338) );
NOR2_X4 U_g27339 ( .A1(g27093), .A2(g26464), .ZN(g27339) );
NOR2_X4 U_g27340 ( .A1(g27096), .A2(g26469), .ZN(g27340) );
NOR2_X4 U_g27341 ( .A1(g27097), .A2(g26470), .ZN(g27341) );
NOR2_X4 U_g27342 ( .A1(g27098), .A2(g26473), .ZN(g27342) );
NOR2_X4 U_g27343 ( .A1(g27099), .A2(g26477), .ZN(g27343) );
NOR2_X4 U_g27344 ( .A1(g27100), .A2(g26478), .ZN(g27344) );
NOR2_X4 U_g27345 ( .A1(g27101), .A2(g26479), .ZN(g27345) );
NOR2_X4 U_g27346 ( .A1(g27105), .A2(g26488), .ZN(g27346) );
NOR2_X4 U_g27347 ( .A1(g27108), .A2(g26493), .ZN(g27347) );
NOR2_X4 U_g27348 ( .A1(g27109), .A2(g26494), .ZN(g27348) );
NOR2_X4 U_g27354 ( .A1(g27112), .A2(g26504), .ZN(g27354) );
NOR2_X4 U_g27414 ( .A1(g26770), .A2(g25187), .ZN(g27414) );
NOR3_X4 U_g27415 ( .A1(g23104), .A2(g27181), .A3(g25128), .ZN(g27415) );
NOR2_X4 U_g27435 ( .A1(g26777), .A2(g25193), .ZN(g27435) );
NOR3_X4 U_g27436 ( .A1(g23118), .A2(g27187), .A3(g24427), .ZN(g27436) );
NOR2_X4 U_g27450 ( .A1(g26902), .A2(g24613), .ZN(g27450) );
NOR2_X4 U_g27454 ( .A1(g26783), .A2(g25196), .ZN(g27454) );
NOR3_X4 U_g27455 ( .A1(g23127), .A2(g26758), .A3(g24431), .ZN(g27455) );
NOR2_X4 U_g27462 ( .A1(g26892), .A2(g24622), .ZN(g27462) );
NOR2_X4 U_g27464 ( .A1(g27178), .A2(g25975), .ZN(g27464) );
NOR2_X4 U_g27466 ( .A1(g26915), .A2(g24624), .ZN(g27466) );
NOR2_X4 U_g27470 ( .A1(g26790), .A2(g25198), .ZN(g27470) );
NOR3_X4 U_g27471 ( .A1(g23138), .A2(g26764), .A3(g24435), .ZN(g27471) );
NOR2_X4 U_g27478 ( .A1(g26754), .A2(g24432), .ZN(g27478) );
NOR2_X4 U_g27481 ( .A1(g27182), .A2(g25980), .ZN(g27481) );
NOR2_X4 U_g27482 ( .A1(g26906), .A2(g24637), .ZN(g27482) );
NOR2_X4 U_g27485 ( .A1(g26928), .A2(g24638), .ZN(g27485) );
NOR3_X4 U_g27492 ( .A1(g24958), .A2(g24633), .A3(g26771), .ZN(g27492) );
NOR2_X4 U_g27496 ( .A1(g27185), .A2(g25178), .ZN(g27496) );
NOR2_X4 U_g27501 ( .A1(g26763), .A2(g24436), .ZN(g27501) );
NOR2_X4 U_g27504 ( .A1(g26918), .A2(g24656), .ZN(g27504) );
NOR2_X4 U_g27507 ( .A1(g26941), .A2(g24657), .ZN(g27507) );
NOR3_X4 U_g27513 ( .A1(g24969), .A2(g24653), .A3(g26778), .ZN(g27513) );
NOR2_X4 U_g27521 ( .A1(g26766), .A2(g24439), .ZN(g27521) );
NOR2_X4 U_g27524 ( .A1(g26931), .A2(g24675), .ZN(g27524) );
NOR2_X4 U_g27527 ( .A1(g26759), .A2(g19087), .ZN(g27527) );
NOR2_X4 U_g27529 ( .A1(g4456), .A2(g26873), .ZN(g27529) );
NOR2_X4 U_g27531 ( .A1(g26760), .A2(g25181), .ZN(g27531) );
NOR2_X4 U_g27532 ( .A1(g26761), .A2(g25182), .ZN(g27532) );
NOR3_X4 U_g27538 ( .A1(g24982), .A2(g24672), .A3(g26784), .ZN(g27538) );
NOR2_X4 U_g27546 ( .A1(g26769), .A2(g24441), .ZN(g27546) );
NOR2_X4 U_g27549 ( .A1(g26765), .A2(g19093), .ZN(g27549) );
NOR2_X4 U_g27551 ( .A1(g4632), .A2(g26882), .ZN(g27551) );
NOR3_X4 U_g27558 ( .A1(g24993), .A2(g24691), .A3(g26791), .ZN(g27558) );
NOR2_X4 U_g27563 ( .A1(g26922), .A2(g24708), .ZN(g27563) );
NOR2_X4 U_g27564 ( .A1(g26767), .A2(g25184), .ZN(g27564) );
NOR2_X4 U_g27565 ( .A1(g26768), .A2(g19100), .ZN(g27565) );
NOR2_X4 U_g27567 ( .A1(g4809), .A2(g26891), .ZN(g27567) );
NOR2_X4 U_g27572 ( .A1(g26911), .A2(g24717), .ZN(g27572) );
NOR2_X4 U_g27573 ( .A1(g26773), .A2(g25188), .ZN(g27573) );
NOR2_X4 U_g27574 ( .A1(g26935), .A2(g24720), .ZN(g27574) );
NOR2_X4 U_g27575 ( .A1(g26774), .A2(g19107), .ZN(g27575) );
NOR2_X4 U_g27577 ( .A1(g4985), .A2(g26901), .ZN(g27577) );
NOR2_X4 U_g27579 ( .A1(g26775), .A2(g25192), .ZN(g27579) );
NOR2_X4 U_g27581 ( .A1(g26925), .A2(g24728), .ZN(g27581) );
NOR2_X4 U_g27582 ( .A1(g26944), .A2(g24731), .ZN(g27582) );
NOR2_X4 U_g27584 ( .A1(g26938), .A2(g24736), .ZN(g27584) );
NOR2_X4 U_g27585 ( .A1(g26950), .A2(g24739), .ZN(g27585) );
NOR2_X4 U_g27588 ( .A1(g26947), .A2(g24742), .ZN(g27588) );
NOR2_X4 U_g27594 ( .A1(g27175), .A2(g17001), .ZN(g27594) );
NOR2_X4 U_g27603 ( .A1(g27179), .A2(g17031), .ZN(g27603) );
NOR2_X4 U_g27612 ( .A1(g27184), .A2(g17065), .ZN(g27612) );
NOR2_X4 U_g27621 ( .A1(g27188), .A2(g17100), .ZN(g27621) );
NOR2_X4 U_g27629 ( .A1(g26829), .A2(g26051), .ZN(g27629) );
NOR2_X4 U_g27631 ( .A1(g26833), .A2(g26053), .ZN(g27631) );
NOR2_X4 U_g27655 ( .A1(g26842), .A2(g26061), .ZN(g27655) );
NOR2_X4 U_g27658 ( .A1(g26851), .A2(g26068), .ZN(g27658) );
NOR2_X4 U_g27672 ( .A1(g26799), .A2(g10024), .ZN(g27672) );
NOR2_X4 U_g27678 ( .A1(g26800), .A2(g10133), .ZN(g27678) );
NOR2_X4 U_g27682 ( .A1(g26801), .A2(g10238), .ZN(g27682) );
NOR2_X4 U_g27718 ( .A1(g27251), .A2(g10133), .ZN(g27718) );
NOR2_X4 U_g27722 ( .A1(g27252), .A2(g10238), .ZN(g27722) );
NOR2_X4 U_g27724 ( .A1(g27254), .A2(g10340), .ZN(g27724) );
NOR2_X4 U_g27735 ( .A1(g27394), .A2(g26961), .ZN(g27735) );
NOR2_X4 U_g27736 ( .A1(g27396), .A2(g26962), .ZN(g27736) );
NOR2_X4 U_g27741 ( .A1(g27407), .A2(g26966), .ZN(g27741) );
NOR2_X4 U_g27742 ( .A1(g27409), .A2(g26967), .ZN(g27742) );
NOR2_X4 U_g27746 ( .A1(g27425), .A2(g26972), .ZN(g27746) );
NOR2_X4 U_g27747 ( .A1(g27427), .A2(g26973), .ZN(g27747) );
NOR2_X4 U_g27754 ( .A1(g27446), .A2(g26985), .ZN(g27754) );
NOR2_X4 U_g27755 ( .A1(g27448), .A2(g26986), .ZN(g27755) );
NOR2_X4 U_g27759 ( .A1(g27495), .A2(g27052), .ZN(g27759) );
NOR2_X4 U_g27760 ( .A1(g27509), .A2(g27076), .ZN(g27760) );
NOR2_X4 U_g27761 ( .A1(g27516), .A2(g27079), .ZN(g27761) );
NOR2_X4 U_g27762 ( .A1(g27530), .A2(g27091), .ZN(g27762) );
NOR2_X4 U_g27763 ( .A1(g27534), .A2(g27092), .ZN(g27763) );
NOR2_X4 U_g27764 ( .A1(g27541), .A2(g27095), .ZN(g27764) );
NOR2_X4 U_g27765 ( .A1(g27552), .A2(g27103), .ZN(g27765) );
NOR2_X4 U_g27766 ( .A1(g27554), .A2(g27104), .ZN(g27766) );
NOR2_X4 U_g27767 ( .A1(g27561), .A2(g27107), .ZN(g27767) );
NOR2_X4 U_g27768 ( .A1(g27568), .A2(g27110), .ZN(g27768) );
NOR2_X4 U_g27769 ( .A1(g27570), .A2(g27111), .ZN(g27769) );
NOR2_X4 U_g27771 ( .A1(g27578), .A2(g27115), .ZN(g27771) );
NOR2_X4 U_g27798 ( .A1(g27632), .A2(g1223), .ZN(g27798) );
NOR3_X4 U_g27802 ( .A1(g6087), .A2(g27632), .A3(g25330), .ZN(g27802) );
NOR2_X4 U_g27810 ( .A1(g27632), .A2(g1215), .ZN(g27810) );
NOR3_X4 U_g27811 ( .A1(g6087), .A2(g27632), .A3(g25404), .ZN(g27811) );
NOR3_X4 U_g27814 ( .A1(g6087), .A2(g27632), .A3(g25322), .ZN(g27814) );
NOR2_X4 U_g27823 ( .A1(g27632), .A2(g1216), .ZN(g27823) );
NOR3_X4 U_g27824 ( .A1(g6087), .A2(g27632), .A3(g25399), .ZN(g27824) );
NOR3_X4 U_g27827 ( .A1(g6087), .A2(g27632), .A3(g25314), .ZN(g27827) );
NOR2_X4 U_g27834 ( .A1(g27478), .A2(g14630), .ZN(g27834) );
NOR2_X4 U_g27842 ( .A1(g27632), .A2(g1217), .ZN(g27842) );
NOR2_X4 U_g27850 ( .A1(g27501), .A2(g14650), .ZN(g27850) );
NOR2_X4 U_g27854 ( .A1(g27632), .A2(g1218), .ZN(g27854) );
NOR3_X4 U_g27855 ( .A1(g6087), .A2(g27632), .A3(g25385), .ZN(g27855) );
NOR2_X4 U_g27864 ( .A1(g27632), .A2(g1219), .ZN(g27864) );
NOR3_X4 U_g27865 ( .A1(g6087), .A2(g27632), .A3(g25370), .ZN(g27865) );
NOR2_X4 U_g27868 ( .A1(g23742), .A2(g27632), .ZN(g27868) );
NOR2_X4 U_g27869 ( .A1(g27632), .A2(g25437), .ZN(g27869) );
NOR2_X4 U_g27875 ( .A1(g27521), .A2(g14677), .ZN(g27875) );
NOR2_X4 U_g27882 ( .A1(g27632), .A2(g1220), .ZN(g27882) );
NOR3_X4 U_g27883 ( .A1(g6087), .A2(g27632), .A3(g25361), .ZN(g27883) );
NOR2_X4 U_g27886 ( .A1(g27632), .A2(g24627), .ZN(g27886) );
NOR2_X4 U_g27892 ( .A1(g27546), .A2(g14711), .ZN(g27892) );
NOR2_X4 U_g27896 ( .A1(g27632), .A2(g1222), .ZN(g27896) );
NOR3_X4 U_g27897 ( .A1(g6087), .A2(g27632), .A3(g25349), .ZN(g27897) );
NOR3_X4 U_g27900 ( .A1(g6087), .A2(g27632), .A3(g25338), .ZN(g27900) );
NOR2_X4 U_g27906 ( .A1(g16127), .A2(g27656), .ZN(g27906) );
NOR2_X4 U_g27911 ( .A1(g16170), .A2(g27657), .ZN(g27911) );
NOR2_X4 U_g27916 ( .A1(g16219), .A2(g27659), .ZN(g27916) );
NOR2_X4 U_g27917 ( .A1(g16220), .A2(g27660), .ZN(g27917) );
NOR2_X4 U_g27925 ( .A1(g16276), .A2(g27661), .ZN(g27925) );
NOR2_X4 U_g27937 ( .A1(g16321), .A2(g27666), .ZN(g27937) );
NOR2_X4 U_g27950 ( .A1(g16367), .A2(g27673), .ZN(g27950) );
NOR2_X4 U_g27962 ( .A1(g16394), .A2(g27679), .ZN(g27962) );
NOR2_X4 U_g27964 ( .A1(g16400), .A2(g27680), .ZN(g27964) );
NOR2_X4 U_g27980 ( .A1(g16428), .A2(g27681), .ZN(g27980) );
NOR2_X4 U_g27997 ( .A1(g16456), .A2(g27242), .ZN(g27997) );
NOR2_X4 U_g28002 ( .A1(g26032), .A2(g27246), .ZN(g28002) );
NOR2_X4 U_g28029 ( .A1(g26033), .A2(g27247), .ZN(g28029) );
NOR2_X4 U_g28059 ( .A1(g26034), .A2(g27248), .ZN(g28059) );
NOR2_X4 U_g28088 ( .A1(g26036), .A2(g27249), .ZN(g28088) );
NOR2_X4 U_g28145 ( .A1(g27629), .A2(g17001), .ZN(g28145) );
NOR2_X4 U_g28146 ( .A1(g27631), .A2(g17031), .ZN(g28146) );
NOR2_X4 U_g28147 ( .A1(g27655), .A2(g17065), .ZN(g28147) );
NOR2_X4 U_g28148 ( .A1(g27658), .A2(g17100), .ZN(g28148) );
NOR2_X4 U_g28157 ( .A1(g13902), .A2(g27370), .ZN(g28157) );
NOR2_X4 U_g28185 ( .A1(g27356), .A2(g26845), .ZN(g28185) );
NOR2_X4 U_g28189 ( .A1(g27359), .A2(g26853), .ZN(g28189) );
NOR2_X4 U_g28191 ( .A1(g27365), .A2(g26860), .ZN(g28191) );
NOR2_X4 U_g28192 ( .A1(g27372), .A2(g26866), .ZN(g28192) );
NOR2_X4 U_g28199 ( .A1(g27250), .A2(g10024), .ZN(g28199) );
NOR2_X4 U_g28321 ( .A1(g27742), .A2(g10133), .ZN(g28321) );
NOR2_X4 U_g28325 ( .A1(g27747), .A2(g10238), .ZN(g28325) );
NOR2_X4 U_g28328 ( .A1(g27755), .A2(g10340), .ZN(g28328) );
NOR2_X4 U_g28342 ( .A1(g15460), .A2(g28008), .ZN(g28342) );
NOR2_X4 U_g28344 ( .A1(g15526), .A2(g28027), .ZN(g28344) );
NOR2_X4 U_g28345 ( .A1(g15527), .A2(g28028), .ZN(g28345) );
NOR2_X4 U_g28346 ( .A1(g15546), .A2(g28035), .ZN(g28346) );
NOR2_X4 U_g28348 ( .A1(g15594), .A2(g28050), .ZN(g28348) );
NOR2_X4 U_g28349 ( .A1(g15595), .A2(g28051), .ZN(g28349) );
NOR2_X4 U_g28350 ( .A1(g15604), .A2(g28057), .ZN(g28350) );
NOR2_X4 U_g28351 ( .A1(g15605), .A2(g28058), .ZN(g28351) );
NOR2_X4 U_g28352 ( .A1(g15624), .A2(g28065), .ZN(g28352) );
NOR2_X4 U_g28353 ( .A1(g15666), .A2(g28073), .ZN(g28353) );
NOR2_X4 U_g28354 ( .A1(g15670), .A2(g28079), .ZN(g28354) );
NOR2_X4 U_g28355 ( .A1(g15671), .A2(g28080), .ZN(g28355) );
NOR2_X4 U_g28356 ( .A1(g15680), .A2(g28086), .ZN(g28356) );
NOR2_X4 U_g28357 ( .A1(g15681), .A2(g28087), .ZN(g28357) );
NOR2_X4 U_g28358 ( .A1(g15700), .A2(g28094), .ZN(g28358) );
NOR2_X4 U_g28360 ( .A1(g15725), .A2(g28098), .ZN(g28360) );
NOR2_X4 U_g28361 ( .A1(g15729), .A2(g28104), .ZN(g28361) );
NOR2_X4 U_g28362 ( .A1(g15730), .A2(g28105), .ZN(g28362) );
NOR2_X4 U_g28363 ( .A1(g15739), .A2(g28111), .ZN(g28363) );
NOR2_X4 U_g28364 ( .A1(g15740), .A2(g28112), .ZN(g28364) );
NOR2_X4 U_g28366 ( .A1(g15765), .A2(g28116), .ZN(g28366) );
NOR2_X4 U_g28367 ( .A1(g15769), .A2(g28122), .ZN(g28367) );
NOR2_X4 U_g28368 ( .A1(g15770), .A2(g28123), .ZN(g28368) );
NOR2_X4 U_g28371 ( .A1(g15793), .A2(g28127), .ZN(g28371) );
NOR2_X4 U_g28392 ( .A1(g27886), .A2(g22344), .ZN(g28392) );
NOR2_X4 U_g28394 ( .A1(g27869), .A2(g22344), .ZN(g28394) );
NOR2_X4 U_g28397 ( .A1(g27869), .A2(g22344), .ZN(g28397) );
NOR2_X4 U_g28400 ( .A1(g27886), .A2(g22344), .ZN(g28400) );
NOR2_X4 U_g28403 ( .A1(g27811), .A2(g22344), .ZN(g28403) );
NOR2_X4 U_g28406 ( .A1(g27824), .A2(g22344), .ZN(g28406) );
NOR2_X4 U_g28409 ( .A1(g24676), .A2(g27801), .ZN(g28409) );
NOR2_X4 U_g28410 ( .A1(g27748), .A2(g22344), .ZN(g28410) );
NOR2_X4 U_g28413 ( .A1(g24695), .A2(g27809), .ZN(g28413) );
NOR2_X4 U_g28414 ( .A1(g27748), .A2(g22344), .ZN(g28414) );
NOR2_X4 U_g28417 ( .A1(g24712), .A2(g27830), .ZN(g28417) );
NOR2_X4 U_g28418 ( .A1(g24723), .A2(g27846), .ZN(g28418) );
NOR2_X4 U_g28420 ( .A1(g16031), .A2(g28171), .ZN(g28420) );
NOR2_X4 U_g28421 ( .A1(g16068), .A2(g28176), .ZN(g28421) );
NOR2_X4 U_g28425 ( .A1(g16133), .A2(g28188), .ZN(g28425) );
NOR2_X4 U_g28449 ( .A1(g27727), .A2(g26780), .ZN(g28449) );
NOR2_X4 U_g28461 ( .A1(g27729), .A2(g26787), .ZN(g28461) );
NOR2_X4 U_g28470 ( .A1(g27671), .A2(g28193), .ZN(g28470) );
NOR2_X4 U_g28473 ( .A1(g27730), .A2(g26794), .ZN(g28473) );
NOR2_X4 U_g28482 ( .A1(g27731), .A2(g26797), .ZN(g28482) );
NOR2_X4 U_g28488 ( .A1(g26755), .A2(g27719), .ZN(g28488) );
NOR2_X4 U_g28489 ( .A1(g26756), .A2(g27720), .ZN(g28489) );
NOR2_X4 U_g28490 ( .A1(g27240), .A2(g27721), .ZN(g28490) );
NOR2_X4 U_g28495 ( .A1(g27244), .A2(g27723), .ZN(g28495) );
NOR2_X4 U_g28499 ( .A1(g26027), .A2(g27725), .ZN(g28499) );
NOR2_X4 U_g28523 ( .A1(g26035), .A2(g27732), .ZN(g28523) );
NOR2_X4 U_g28525 ( .A1(g27245), .A2(g27726), .ZN(g28525) );
NOR2_X4 U_g28528 ( .A1(g26030), .A2(g27728), .ZN(g28528) );
NOR2_X4 U_g28551 ( .A1(g26038), .A2(g27733), .ZN(g28551) );
NOR2_X4 U_g28578 ( .A1(g26039), .A2(g27734), .ZN(g28578) );
NOR2_X4 U_g28606 ( .A1(g26040), .A2(g27737), .ZN(g28606) );
NOR2_X4 U_g28634 ( .A1(g28185), .A2(g17001), .ZN(g28634) );
NOR2_X4 U_g28635 ( .A1(g28189), .A2(g17031), .ZN(g28635) );
NOR2_X4 U_g28636 ( .A1(g28191), .A2(g17065), .ZN(g28636) );
NOR2_X4 U_g28637 ( .A1(g28192), .A2(g17100), .ZN(g28637) );
NOR2_X4 U_g28654 ( .A1(g27770), .A2(g27355), .ZN(g28654) );
NOR2_X4 U_g28656 ( .A1(g27772), .A2(g27358), .ZN(g28656) );
NOR2_X4 U_g28658 ( .A1(g27773), .A2(g27364), .ZN(g28658) );
NOR2_X4 U_g28661 ( .A1(g27775), .A2(g27371), .ZN(g28661) );
NOR2_X4 U_g28668 ( .A1(g27736), .A2(g10024), .ZN(g28668) );
NOR2_X4 U_g28728 ( .A1(g28422), .A2(g27904), .ZN(g28728) );
NOR2_X4 U_g28731 ( .A1(g28423), .A2(g27908), .ZN(g28731) );
NOR2_X4 U_g28732 ( .A1(g14894), .A2(g28426), .ZN(g28732) );
NOR2_X4 U_g28733 ( .A1(g28424), .A2(g27909), .ZN(g28733) );
NOR2_X4 U_g28735 ( .A1(g14957), .A2(g28430), .ZN(g28735) );
NOR2_X4 U_g28736 ( .A1(g28427), .A2(g27913), .ZN(g28736) );
NOR2_X4 U_g28737 ( .A1(g28428), .A2(g27914), .ZN(g28737) );
NOR2_X4 U_g28738 ( .A1(g14975), .A2(g28433), .ZN(g28738) );
NOR2_X4 U_g28739 ( .A1(g28429), .A2(g27915), .ZN(g28739) );
NOR2_X4 U_g28744 ( .A1(g15030), .A2(g28439), .ZN(g28744) );
NOR2_X4 U_g28745 ( .A1(g28431), .A2(g27922), .ZN(g28745) );
NOR2_X4 U_g28746 ( .A1(g15046), .A2(g28441), .ZN(g28746) );
NOR2_X4 U_g28747 ( .A1(g28434), .A2(g27923), .ZN(g28747) );
NOR2_X4 U_g28748 ( .A1(g28435), .A2(g27924), .ZN(g28748) );
NOR2_X4 U_g28749 ( .A1(g15064), .A2(g28444), .ZN(g28749) );
NOR2_X4 U_g28750 ( .A1(g28436), .A2(g27926), .ZN(g28750) );
NOR2_X4 U_g28754 ( .A1(g28440), .A2(g27931), .ZN(g28754) );
NOR2_X4 U_g28758 ( .A1(g15126), .A2(g28451), .ZN(g28758) );
NOR2_X4 U_g28759 ( .A1(g28442), .A2(g27935), .ZN(g28759) );
NOR2_X4 U_g28760 ( .A1(g15142), .A2(g28453), .ZN(g28760) );
NOR2_X4 U_g28761 ( .A1(g28445), .A2(g27936), .ZN(g28761) );
NOR2_X4 U_g28762 ( .A1(g28446), .A2(g27938), .ZN(g28762) );
NOR2_X4 U_g28763 ( .A1(g15160), .A2(g28456), .ZN(g28763) );
NOR2_X4 U_g28767 ( .A1(g28452), .A2(g27945), .ZN(g28767) );
NOR2_X4 U_g28771 ( .A1(g15218), .A2(g28463), .ZN(g28771) );
NOR2_X4 U_g28772 ( .A1(g28454), .A2(g27949), .ZN(g28772) );
NOR2_X4 U_g28773 ( .A1(g15234), .A2(g28465), .ZN(g28773) );
NOR2_X4 U_g28774 ( .A1(g28457), .A2(g27951), .ZN(g28774) );
NOR2_X4 U_g28778 ( .A1(g28464), .A2(g27963), .ZN(g28778) );
NOR2_X4 U_g28782 ( .A1(g15304), .A2(g28475), .ZN(g28782) );
NOR2_X4 U_g28783 ( .A1(g28466), .A2(g27968), .ZN(g28783) );
NOR2_X4 U_g28784 ( .A1(g28468), .A2(g27970), .ZN(g28784) );
NOR2_X4 U_g28788 ( .A1(g28476), .A2(g27984), .ZN(g28788) );
NOR2_X4 U_g28789 ( .A1(g28477), .A2(g27985), .ZN(g28789) );
NOR2_X4 U_g28790 ( .A1(g28478), .A2(g27991), .ZN(g28790) );
NOR2_X4 U_g28794 ( .A1(g28484), .A2(g28009), .ZN(g28794) );
NOR2_X4 U_g28795 ( .A1(g28485), .A2(g28015), .ZN(g28795) );
NOR2_X4 U_g28802 ( .A1(g28492), .A2(g28036), .ZN(g28802) );
NOR2_X4 U_g28803 ( .A1(g28493), .A2(g28042), .ZN(g28803) );
NOR2_X4 U_g28813 ( .A1(g28497), .A2(g28066), .ZN(g28813) );
NOR2_X4 U_g28874 ( .A1(g28657), .A2(g16221), .ZN(g28874) );
NOR2_X4 U_g28886 ( .A1(g28659), .A2(g16277), .ZN(g28886) );
NOR2_X4 U_g28903 ( .A1(g28660), .A2(g13295), .ZN(g28903) );
NOR2_X4 U_g28920 ( .A1(g28662), .A2(g13322), .ZN(g28920) );
NOR2_X4 U_g28941 ( .A1(g28663), .A2(g13343), .ZN(g28941) );
NOR3_X4 U_g28954 ( .A1(g26673), .A2(g27241), .A3(g28323), .ZN(g28954) );
NOR2_X4 U_g28963 ( .A1(g28664), .A2(g13365), .ZN(g28963) );
NOR2_X4 U_g28982 ( .A1(g28665), .A2(g28670), .ZN(g28982) );
NOR2_X4 U_g28987 ( .A1(g28666), .A2(g13390), .ZN(g28987) );
NOR2_X4 U_g28990 ( .A1(g28667), .A2(g16457), .ZN(g28990) );
NOR2_X4 U_g29009 ( .A1(g28669), .A2(g28320), .ZN(g29009) );
NOR2_X4 U_g29013 ( .A1(g28671), .A2(g11607), .ZN(g29013) );
NOR2_X4 U_g29016 ( .A1(g28672), .A2(g13487), .ZN(g29016) );
NOR2_X4 U_g29031 ( .A1(g28319), .A2(g28324), .ZN(g29031) );
NOR2_X4 U_g29039 ( .A1(g28322), .A2(g13500), .ZN(g29039) );
NOR2_X4 U_g29063 ( .A1(g28326), .A2(g28329), .ZN(g29063) );
NOR2_X4 U_g29064 ( .A1(g28327), .A2(g28330), .ZN(g29064) );
NOR2_X4 U_g29083 ( .A1(g28331), .A2(g28333), .ZN(g29083) );
NOR2_X4 U_g29090 ( .A1(g28332), .A2(g28334), .ZN(g29090) );
NOR2_X4 U_g29097 ( .A1(g28335), .A2(g28336), .ZN(g29097) );
NOR2_X4 U_g29109 ( .A1(g28654), .A2(g17001), .ZN(g29109) );
NOR2_X4 U_g29110 ( .A1(g28656), .A2(g17031), .ZN(g29110) );
NOR2_X4 U_g29111 ( .A1(g28658), .A2(g17065), .ZN(g29111) );
NOR2_X4 U_g29112 ( .A1(g28661), .A2(g17100), .ZN(g29112) );
NOR2_X4 U_g29113 ( .A1(g28381), .A2(g8907), .ZN(g29113) );
NOR2_X4 U_g29126 ( .A1(g28373), .A2(g27774), .ZN(g29126) );
NOR2_X4 U_g29127 ( .A1(g28376), .A2(g27779), .ZN(g29127) );
NOR2_X4 U_g29128 ( .A1(g28380), .A2(g27783), .ZN(g29128) );
NOR2_X4 U_g29129 ( .A1(g28385), .A2(g27790), .ZN(g29129) );
NOR2_X4 U_g29167 ( .A1(g28841), .A2(g28396), .ZN(g29167) );
NOR2_X4 U_g29169 ( .A1(g28843), .A2(g28398), .ZN(g29169) );
NOR2_X4 U_g29170 ( .A1(g28844), .A2(g28399), .ZN(g29170) );
NOR2_X4 U_g29172 ( .A1(g28846), .A2(g28401), .ZN(g29172) );
NOR2_X4 U_g29173 ( .A1(g28847), .A2(g28402), .ZN(g29173) );
NOR2_X4 U_g29178 ( .A1(g28848), .A2(g28404), .ZN(g29178) );
NOR2_X4 U_g29179 ( .A1(g28849), .A2(g28405), .ZN(g29179) );
NOR2_X4 U_g29181 ( .A1(g28850), .A2(g28407), .ZN(g29181) );
NOR2_X4 U_g29182 ( .A1(g28851), .A2(g28408), .ZN(g29182) );
NOR2_X4 U_g29184 ( .A1(g28852), .A2(g28411), .ZN(g29184) );
NOR2_X4 U_g29185 ( .A1(g28853), .A2(g28412), .ZN(g29185) );
NOR2_X4 U_g29187 ( .A1(g28854), .A2(g28416), .ZN(g29187) );
NOR2_X4 U_g29194 ( .A1(g14958), .A2(g28881), .ZN(g29194) );
NOR2_X4 U_g29195 ( .A1(g28880), .A2(g28438), .ZN(g29195) );
NOR2_X4 U_g29197 ( .A1(g15031), .A2(g28893), .ZN(g29197) );
NOR2_X4 U_g29198 ( .A1(g15047), .A2(g28898), .ZN(g29198) );
NOR2_X4 U_g29199 ( .A1(g28892), .A2(g28448), .ZN(g29199) );
NOR2_X4 U_g29201 ( .A1(g15104), .A2(g28910), .ZN(g29201) );
NOR2_X4 U_g29202 ( .A1(g28897), .A2(g28450), .ZN(g29202) );
NOR2_X4 U_g29204 ( .A1(g15127), .A2(g28915), .ZN(g29204) );
NOR2_X4 U_g29205 ( .A1(g15143), .A2(g28923), .ZN(g29205) );
NOR2_X4 U_g29206 ( .A1(g28909), .A2(g28459), .ZN(g29206) );
NOR2_X4 U_g29207 ( .A1(g28914), .A2(g28460), .ZN(g29207) );
NOR2_X4 U_g29209 ( .A1(g15196), .A2(g28936), .ZN(g29209) );
NOR2_X4 U_g29210 ( .A1(g28919), .A2(g28462), .ZN(g29210) );
NOR2_X4 U_g29212 ( .A1(g15219), .A2(g28944), .ZN(g29212) );
NOR2_X4 U_g29213 ( .A1(g15235), .A2(g28949), .ZN(g29213) );
NOR2_X4 U_g29214 ( .A1(g28931), .A2(g28469), .ZN(g29214) );
NOR2_X4 U_g29215 ( .A1(g28935), .A2(g28471), .ZN(g29215) );
NOR2_X4 U_g29216 ( .A1(g28940), .A2(g28472), .ZN(g29216) );
NOR2_X4 U_g29218 ( .A1(g15282), .A2(g28966), .ZN(g29218) );
NOR2_X4 U_g29219 ( .A1(g28948), .A2(g28474), .ZN(g29219) );
NOR2_X4 U_g29221 ( .A1(g15305), .A2(g28971), .ZN(g29221) );
NOR2_X4 U_g29222 ( .A1(g28958), .A2(g28479), .ZN(g29222) );
NOR2_X4 U_g29223 ( .A1(g28962), .A2(g28480), .ZN(g29223) );
NOR2_X4 U_g29224 ( .A1(g28970), .A2(g28481), .ZN(g29224) );
NOR2_X4 U_g29226 ( .A1(g15374), .A2(g28997), .ZN(g29226) );
NOR2_X4 U_g29227 ( .A1(g28986), .A2(g28486), .ZN(g29227) );
NOR2_X4 U_g29228 ( .A1(g28996), .A2(g28487), .ZN(g29228) );
NOR2_X4 U_g29231 ( .A1(g29022), .A2(g28494), .ZN(g29231) );
NOR2_X4 U_g29303 ( .A1(g28716), .A2(g19112), .ZN(g29303) );
NOR2_X4 U_g29313 ( .A1(g28717), .A2(g19117), .ZN(g29313) );
NOR2_X4 U_g29324 ( .A1(g28718), .A2(g19124), .ZN(g29324) );
NOR2_X4 U_g29333 ( .A1(g28719), .A2(g19131), .ZN(g29333) );
NOR2_X4 U_g29340 ( .A1(g28337), .A2(g28722), .ZN(g29340) );
NOR2_X4 U_g29343 ( .A1(g28338), .A2(g28724), .ZN(g29343) );
NOR2_X4 U_g29345 ( .A1(g28339), .A2(g28726), .ZN(g29345) );
NOR2_X4 U_g29347 ( .A1(g28340), .A2(g28729), .ZN(g29347) );
NOR2_X4 U_g29353 ( .A1(g29126), .A2(g17001), .ZN(g29353) );
NOR2_X4 U_g29354 ( .A1(g29127), .A2(g17031), .ZN(g29354) );
NOR2_X4 U_g29355 ( .A1(g29128), .A2(g17065), .ZN(g29355) );
NOR2_X4 U_g29357 ( .A1(g29129), .A2(g17100), .ZN(g29357) );
NOR2_X4 U_g29399 ( .A1(g28834), .A2(g28378), .ZN(g29399) );
NOR2_X4 U_g29403 ( .A1(g28836), .A2(g28383), .ZN(g29403) );
NOR2_X4 U_g29406 ( .A1(g28838), .A2(g28387), .ZN(g29406) );
NOR2_X4 U_g29409 ( .A1(g28840), .A2(g28389), .ZN(g29409) );
NOR2_X4 U_g29552 ( .A1(g29130), .A2(g29411), .ZN(g29552) );
NOR2_X4 U_g29569 ( .A1(g28708), .A2(g29174), .ZN(g29569) );
NOR2_X4 U_g29570 ( .A1(g28709), .A2(g29175), .ZN(g29570) );
NOR2_X4 U_g29571 ( .A1(g28710), .A2(g29176), .ZN(g29571) );
NOR2_X4 U_g29574 ( .A1(g28712), .A2(g29180), .ZN(g29574) );
NOR2_X4 U_g29576 ( .A1(g28713), .A2(g29183), .ZN(g29576) );
NOR2_X4 U_g29577 ( .A1(g28714), .A2(g29186), .ZN(g29577) );
NOR2_X4 U_g29578 ( .A1(g28715), .A2(g29188), .ZN(g29578) );
NOR2_X4 U_g29579 ( .A1(g29399), .A2(g17001), .ZN(g29579) );
NOR2_X4 U_g29580 ( .A1(g29403), .A2(g17031), .ZN(g29580) );
NOR2_X4 U_g29581 ( .A1(g29406), .A2(g17065), .ZN(g29581) );
NOR2_X4 U_g29582 ( .A1(g29409), .A2(g17100), .ZN(g29582) );
NOR2_X4 U_g29606 ( .A1(g13878), .A2(g29248), .ZN(g29606) );
NOR2_X4 U_g29608 ( .A1(g13892), .A2(g29251), .ZN(g29608) );
NOR2_X4 U_g29609 ( .A1(g13900), .A2(g29252), .ZN(g29609) );
NOR2_X4 U_g29611 ( .A1(g13913), .A2(g29255), .ZN(g29611) );
NOR2_X4 U_g29612 ( .A1(g13933), .A2(g29256), .ZN(g29612) );
NOR2_X4 U_g29613 ( .A1(g13941), .A2(g29257), .ZN(g29613) );
NOR2_X4 U_g29616 ( .A1(g13969), .A2(g29259), .ZN(g29616) );
NOR2_X4 U_g29617 ( .A1(g13989), .A2(g29260), .ZN(g29617) );
NOR2_X4 U_g29618 ( .A1(g13997), .A2(g29261), .ZN(g29618) );
NOR2_X4 U_g29620 ( .A1(g14039), .A2(g29262), .ZN(g29620) );
NOR2_X4 U_g29621 ( .A1(g14059), .A2(g29263), .ZN(g29621) );
NOR2_X4 U_g29623 ( .A1(g14130), .A2(g29264), .ZN(g29623) );
NOR2_X4 U_g29663 ( .A1(g29518), .A2(g29284), .ZN(g29663) );
NOR2_X4 U_g29665 ( .A1(g29521), .A2(g29289), .ZN(g29665) );
NOR2_X4 U_g29667 ( .A1(g29524), .A2(g29294), .ZN(g29667) );
NOR2_X4 U_g29669 ( .A1(g29528), .A2(g29300), .ZN(g29669) );
NOR2_X4 U_g29670 ( .A1(g29529), .A2(g29302), .ZN(g29670) );
NOR2_X4 U_g29671 ( .A1(g29534), .A2(g29310), .ZN(g29671) );
NOR2_X4 U_g29672 ( .A1(g29536), .A2(g29312), .ZN(g29672) );
NOR2_X4 U_g29676 ( .A1(g29540), .A2(g29320), .ZN(g29676) );
NOR2_X4 U_g29677 ( .A1(g29543), .A2(g29321), .ZN(g29677) );
NOR2_X4 U_g29678 ( .A1(g29545), .A2(g29323), .ZN(g29678) );
NOR2_X4 U_g29679 ( .A1(g29549), .A2(g29329), .ZN(g29679) );
NOR2_X4 U_g29680 ( .A1(g29553), .A2(g29330), .ZN(g29680) );
NOR2_X4 U_g29681 ( .A1(g29555), .A2(g29332), .ZN(g29681) );
NOR2_X4 U_g29682 ( .A1(g29557), .A2(g29336), .ZN(g29682) );
NOR2_X4 U_g29683 ( .A1(g29559), .A2(g29337), .ZN(g29683) );
NOR2_X4 U_g29684 ( .A1(g29562), .A2(g29338), .ZN(g29684) );
NOR2_X4 U_g29685 ( .A1(g29564), .A2(g29341), .ZN(g29685) );
NOR2_X4 U_g29686 ( .A1(g29566), .A2(g29342), .ZN(g29686) );
NOR2_X4 U_g29687 ( .A1(g29572), .A2(g29344), .ZN(g29687) );
NOR2_X4 U_g29688 ( .A1(g29575), .A2(g29346), .ZN(g29688) );
NOR2_X4 U_g29703 ( .A1(g29583), .A2(g1917), .ZN(g29703) );
NOR3_X4 U_g29705 ( .A1(g6104), .A2(g29583), .A3(g25339), .ZN(g29705) );
NOR2_X4 U_g29709 ( .A1(g29583), .A2(g1909), .ZN(g29709) );
NOR3_X4 U_g29710 ( .A1(g6104), .A2(g29583), .A3(g25412), .ZN(g29710) );
NOR3_X4 U_g29713 ( .A1(g6104), .A2(g29583), .A3(g25332), .ZN(g29713) );
NOR2_X4 U_g29717 ( .A1(g29583), .A2(g1910), .ZN(g29717) );
NOR3_X4 U_g29718 ( .A1(g6104), .A2(g29583), .A3(g25409), .ZN(g29718) );
NOR3_X4 U_g29721 ( .A1(g6104), .A2(g29583), .A3(g25323), .ZN(g29721) );
NOR2_X4 U_g29725 ( .A1(g29583), .A2(g1911), .ZN(g29725) );
NOR2_X4 U_g29727 ( .A1(g29583), .A2(g1912), .ZN(g29727) );
NOR3_X4 U_g29728 ( .A1(g6104), .A2(g29583), .A3(g25401), .ZN(g29728) );
NOR2_X4 U_g29731 ( .A1(g29583), .A2(g1913), .ZN(g29731) );
NOR3_X4 U_g29732 ( .A1(g6104), .A2(g29583), .A3(g25387), .ZN(g29732) );
NOR2_X4 U_g29735 ( .A1(g23797), .A2(g29583), .ZN(g29735) );
NOR2_X4 U_g29736 ( .A1(g29583), .A2(g25444), .ZN(g29736) );
NOR2_X4 U_g29740 ( .A1(g29583), .A2(g1914), .ZN(g29740) );
NOR3_X4 U_g29741 ( .A1(g6104), .A2(g29583), .A3(g25376), .ZN(g29741) );
NOR2_X4 U_g29744 ( .A1(g29583), .A2(g24641), .ZN(g29744) );
NOR2_X4 U_g29747 ( .A1(g29583), .A2(g1916), .ZN(g29747) );
NOR3_X4 U_g29748 ( .A1(g6104), .A2(g29583), .A3(g25363), .ZN(g29748) );
NOR3_X4 U_g29751 ( .A1(g6104), .A2(g29583), .A3(g25352), .ZN(g29751) );
NOR2_X4 U_g29754 ( .A1(g16178), .A2(g29607), .ZN(g29754) );
NOR2_X4 U_g29755 ( .A1(g16229), .A2(g29610), .ZN(g29755) );
NOR2_X4 U_g29756 ( .A1(g16284), .A2(g29614), .ZN(g29756) );
NOR2_X4 U_g29757 ( .A1(g16285), .A2(g29615), .ZN(g29757) );
NOR2_X4 U_g29758 ( .A1(g16335), .A2(g29619), .ZN(g29758) );
NOR2_X4 U_g29759 ( .A1(g16379), .A2(g29622), .ZN(g29759) );
NOR2_X4 U_g29760 ( .A1(g16411), .A2(g29624), .ZN(g29760) );
NOR3_X4 U_g29761 ( .A1(g28707), .A2(g28711), .A3(g29466), .ZN(g29761) );
NOR2_X4 U_g29762 ( .A1(g16432), .A2(g29625), .ZN(g29762) );
NOR2_X4 U_g29763 ( .A1(g16438), .A2(g29626), .ZN(g29763) );
NOR2_X4 U_g29764 ( .A1(g16462), .A2(g29464), .ZN(g29764) );
NOR2_X4 U_g29765 ( .A1(g13492), .A2(g29465), .ZN(g29765) );
NOR2_X4 U_g29766 ( .A1(g29467), .A2(g19142), .ZN(g29766) );
NOR2_X4 U_g29767 ( .A1(g29468), .A2(g19143), .ZN(g29767) );
NOR2_X4 U_g29768 ( .A1(g29469), .A2(g19146), .ZN(g29768) );
NOR2_X4 U_g29769 ( .A1(g29470), .A2(g19148), .ZN(g29769) );
NOR2_X4 U_g29770 ( .A1(g29471), .A2(g29196), .ZN(g29770) );
NOR2_X4 U_g29771 ( .A1(g29472), .A2(g29200), .ZN(g29771) );
NOR2_X4 U_g29772 ( .A1(g29473), .A2(g29203), .ZN(g29772) );
NOR2_X4 U_g29773 ( .A1(g29474), .A2(g29208), .ZN(g29773) );
NOR2_X4 U_g29774 ( .A1(g29475), .A2(g29211), .ZN(g29774) );
NOR2_X4 U_g29775 ( .A1(g29476), .A2(g29217), .ZN(g29775) );
NOR2_X4 U_g29776 ( .A1(g29477), .A2(g29220), .ZN(g29776) );
NOR2_X4 U_g29777 ( .A1(g29478), .A2(g29225), .ZN(g29777) );
NOR2_X4 U_g29778 ( .A1(g29479), .A2(g29229), .ZN(g29778) );
NOR2_X4 U_g29779 ( .A1(g13943), .A2(g29502), .ZN(g29779) );
NOR2_X4 U_g29780 ( .A1(g29480), .A2(g29232), .ZN(g29780) );
NOR2_X4 U_g29781 ( .A1(g29481), .A2(g29233), .ZN(g29781) );
NOR2_X4 U_g29782 ( .A1(g29482), .A2(g29234), .ZN(g29782) );
NOR2_X4 U_g29783 ( .A1(g29483), .A2(g29235), .ZN(g29783) );
NOR2_X4 U_g29784 ( .A1(g29484), .A2(g29236), .ZN(g29784) );
NOR2_X4 U_g29785 ( .A1(g29485), .A2(g29238), .ZN(g29785) );
NOR2_X4 U_g29786 ( .A1(g29486), .A2(g29239), .ZN(g29786) );
NOR2_X4 U_g29787 ( .A1(g29487), .A2(g29240), .ZN(g29787) );
NOR2_X4 U_g29788 ( .A1(g29488), .A2(g29241), .ZN(g29788) );
NOR2_X4 U_g29789 ( .A1(g29489), .A2(g29242), .ZN(g29789) );
NOR2_X4 U_g29791 ( .A1(g29490), .A2(g29243), .ZN(g29791) );
NOR2_X4 U_g29912 ( .A1(g24676), .A2(g29716), .ZN(g29912) );
NOR2_X4 U_g29914 ( .A1(g24695), .A2(g29724), .ZN(g29914) );
NOR2_X4 U_g29916 ( .A1(g24712), .A2(g29726), .ZN(g29916) );
NOR2_X4 U_g29918 ( .A1(g29744), .A2(g22367), .ZN(g29918) );
NOR2_X4 U_g29919 ( .A1(g29736), .A2(g22367), .ZN(g29919) );
NOR2_X4 U_g29920 ( .A1(g24723), .A2(g29739), .ZN(g29920) );
NOR2_X4 U_g29921 ( .A1(g29736), .A2(g22367), .ZN(g29921) );
NOR2_X4 U_g29922 ( .A1(g29744), .A2(g22367), .ZN(g29922) );
NOR2_X4 U_g29924 ( .A1(g29710), .A2(g22367), .ZN(g29924) );
NOR2_X4 U_g29926 ( .A1(g29718), .A2(g22367), .ZN(g29926) );
NOR2_X4 U_g29928 ( .A1(g29673), .A2(g22367), .ZN(g29928) );
NOR2_X4 U_g29929 ( .A1(g29673), .A2(g22367), .ZN(g29929) );
NOR2_X4 U_g29936 ( .A1(g16049), .A2(g29790), .ZN(g29936) );
NOR2_X4 U_g29939 ( .A1(g16102), .A2(g29792), .ZN(g29939) );
NOR2_X4 U_g29941 ( .A1(g16182), .A2(g29793), .ZN(g29941) );
NOR2_X4 U_g30010 ( .A1(g29520), .A2(g29942), .ZN(g30010) );
NOR2_X4 U_g30011 ( .A1(g29522), .A2(g29944), .ZN(g30011) );
NOR2_X4 U_g30012 ( .A1(g29523), .A2(g29945), .ZN(g30012) );
NOR2_X4 U_g30013 ( .A1(g29525), .A2(g29946), .ZN(g30013) );
NOR2_X4 U_g30014 ( .A1(g29526), .A2(g29947), .ZN(g30014) );
NOR2_X4 U_g30015 ( .A1(g29527), .A2(g29948), .ZN(g30015) );
NOR2_X4 U_g30016 ( .A1(g29531), .A2(g29949), .ZN(g30016) );
NOR2_X4 U_g30017 ( .A1(g29532), .A2(g29950), .ZN(g30017) );
NOR2_X4 U_g30018 ( .A1(g29533), .A2(g29951), .ZN(g30018) );
NOR2_X4 U_g30019 ( .A1(g29538), .A2(g29952), .ZN(g30019) );
NOR2_X4 U_g30020 ( .A1(g29539), .A2(g29953), .ZN(g30020) );
NOR2_X4 U_g30021 ( .A1(g29541), .A2(g29954), .ZN(g30021) );
NOR2_X4 U_g30022 ( .A1(g29547), .A2(g29955), .ZN(g30022) );
NOR2_X4 U_g30023 ( .A1(g29548), .A2(g29956), .ZN(g30023) );
NOR2_X4 U_g30024 ( .A1(g29550), .A2(g29957), .ZN(g30024) );
NOR2_X4 U_g30025 ( .A1(g29558), .A2(g29958), .ZN(g30025) );
NOR2_X4 U_g30026 ( .A1(g29560), .A2(g29959), .ZN(g30026) );
NOR2_X4 U_g30027 ( .A1(g29565), .A2(g29960), .ZN(g30027) );
NOR2_X4 U_g30028 ( .A1(g29567), .A2(g29961), .ZN(g30028) );
NOR2_X4 U_g30029 ( .A1(g29573), .A2(g29962), .ZN(g30029) );
NOR2_X4 U_g30030 ( .A1(g24676), .A2(g29923), .ZN(g30030) );
NOR2_X4 U_g30031 ( .A1(g24695), .A2(g29925), .ZN(g30031) );
NOR2_X4 U_g30032 ( .A1(g24712), .A2(g29927), .ZN(g30032) );
NOR2_X4 U_g30033 ( .A1(g24723), .A2(g29931), .ZN(g30033) );
NOR2_X4 U_g30053 ( .A1(g29963), .A2(g16286), .ZN(g30053) );
NOR2_X4 U_g30054 ( .A1(g29964), .A2(g16336), .ZN(g30054) );
NOR2_X4 U_g30055 ( .A1(g29965), .A2(g13326), .ZN(g30055) );
NOR2_X4 U_g30056 ( .A1(g29966), .A2(g13345), .ZN(g30056) );
NOR2_X4 U_g30057 ( .A1(g29967), .A2(g13368), .ZN(g30057) );
NOR2_X4 U_g30058 ( .A1(g29968), .A2(g13395), .ZN(g30058) );
NOR2_X4 U_g30059 ( .A1(g29969), .A2(g29811), .ZN(g30059) );
NOR2_X4 U_g30060 ( .A1(g29970), .A2(g11612), .ZN(g30060) );
NOR2_X4 U_g30061 ( .A1(g29971), .A2(g13493), .ZN(g30061) );
NOR2_X4 U_g30062 ( .A1(g29810), .A2(g29815), .ZN(g30062) );
NOR2_X4 U_g30063 ( .A1(g29812), .A2(g11637), .ZN(g30063) );
NOR2_X4 U_g30064 ( .A1(g29813), .A2(g13506), .ZN(g30064) );
NOR2_X4 U_g30065 ( .A1(g29814), .A2(g29817), .ZN(g30065) );
NOR2_X4 U_g30066 ( .A1(g29816), .A2(g13517), .ZN(g30066) );
NOR2_X4 U_g30067 ( .A1(g29818), .A2(g29820), .ZN(g30067) );
NOR2_X4 U_g30068 ( .A1(g29819), .A2(g29821), .ZN(g30068) );
NOR2_X4 U_g30069 ( .A1(g29822), .A2(g29828), .ZN(g30069) );
NOR2_X4 U_g30070 ( .A1(g29827), .A2(g29833), .ZN(g30070) );
NOR2_X4 U_g30071 ( .A1(g29834), .A2(g29839), .ZN(g30071) );
NOR2_X4 U_g30072 ( .A1(g29910), .A2(g8947), .ZN(g30072) );
NOR2_X4 U_g30245 ( .A1(g16074), .A2(g30077), .ZN(g30245) );
NOR2_X4 U_g30246 ( .A1(g16107), .A2(g30079), .ZN(g30246) );
NOR2_X4 U_g30247 ( .A1(g16112), .A2(g30080), .ZN(g30247) );
NOR2_X4 U_g30248 ( .A1(g16139), .A2(g30081), .ZN(g30248) );
NOR2_X4 U_g30249 ( .A1(g16158), .A2(g30082), .ZN(g30249) );
NOR2_X4 U_g30250 ( .A1(g16163), .A2(g30083), .ZN(g30250) );
NOR2_X4 U_g30251 ( .A1(g16198), .A2(g30085), .ZN(g30251) );
NOR2_X4 U_g30252 ( .A1(g16217), .A2(g30086), .ZN(g30252) );
NOR2_X4 U_g30253 ( .A1(g16222), .A2(g30087), .ZN(g30253) );
NOR2_X4 U_g30254 ( .A1(g16242), .A2(g30088), .ZN(g30254) );
NOR2_X4 U_g30255 ( .A1(g16263), .A2(g30089), .ZN(g30255) );
NOR2_X4 U_g30256 ( .A1(g16282), .A2(g30090), .ZN(g30256) );
NOR2_X4 U_g30257 ( .A1(g16290), .A2(g30091), .ZN(g30257) );
NOR2_X4 U_g30258 ( .A1(g16291), .A2(g30092), .ZN(g30258) );
NOR2_X4 U_g30259 ( .A1(g16301), .A2(g30093), .ZN(g30259) );
NOR2_X4 U_g30260 ( .A1(g16322), .A2(g30094), .ZN(g30260) );
NOR2_X4 U_g30261 ( .A1(g16342), .A2(g30095), .ZN(g30261) );
NOR2_X4 U_g30262 ( .A1(g16343), .A2(g30096), .ZN(g30262) );
NOR2_X4 U_g30263 ( .A1(g16344), .A2(g30097), .ZN(g30263) );
NOR2_X4 U_g30264 ( .A1(g16348), .A2(g30098), .ZN(g30264) );
NOR2_X4 U_g30265 ( .A1(g16349), .A2(g30099), .ZN(g30265) );
NOR2_X4 U_g30266 ( .A1(g16359), .A2(g30100), .ZN(g30266) );
NOR2_X4 U_g30267 ( .A1(g16380), .A2(g30101), .ZN(g30267) );
NOR2_X4 U_g30268 ( .A1(g16382), .A2(g30102), .ZN(g30268) );
NOR2_X4 U_g30269 ( .A1(g16386), .A2(g30103), .ZN(g30269) );
NOR2_X4 U_g30270 ( .A1(g16387), .A2(g30104), .ZN(g30270) );
NOR2_X4 U_g30271 ( .A1(g16388), .A2(g30105), .ZN(g30271) );
NOR2_X4 U_g30272 ( .A1(g16392), .A2(g30106), .ZN(g30272) );
NOR2_X4 U_g30273 ( .A1(g16393), .A2(g30107), .ZN(g30273) );
NOR2_X4 U_g30274 ( .A1(g16403), .A2(g30108), .ZN(g30274) );
NOR2_X4 U_g30275 ( .A1(g16413), .A2(g30109), .ZN(g30275) );
NOR2_X4 U_g30276 ( .A1(g16415), .A2(g30110), .ZN(g30276) );
NOR2_X4 U_g30277 ( .A1(g16418), .A2(g30111), .ZN(g30277) );
NOR2_X4 U_g30278 ( .A1(g16420), .A2(g30112), .ZN(g30278) );
NOR2_X4 U_g30279 ( .A1(g16424), .A2(g30113), .ZN(g30279) );
NOR2_X4 U_g30280 ( .A1(g16425), .A2(g30114), .ZN(g30280) );
NOR2_X4 U_g30281 ( .A1(g16426), .A2(g30115), .ZN(g30281) );
NOR2_X4 U_g30282 ( .A1(g16430), .A2(g30117), .ZN(g30282) );
NOR2_X4 U_g30283 ( .A1(g16431), .A2(g30118), .ZN(g30283) );
NOR2_X4 U_g30284 ( .A1(g16444), .A2(g29980), .ZN(g30284) );
NOR2_X4 U_g30285 ( .A1(g16447), .A2(g29981), .ZN(g30285) );
NOR2_X4 U_g30286 ( .A1(g16449), .A2(g29982), .ZN(g30286) );
NOR2_X4 U_g30287 ( .A1(g16452), .A2(g29983), .ZN(g30287) );
NOR2_X4 U_g30288 ( .A1(g16454), .A2(g29984), .ZN(g30288) );
NOR2_X4 U_g30289 ( .A1(g16458), .A2(g29985), .ZN(g30289) );
NOR2_X4 U_g30290 ( .A1(g16459), .A2(g29986), .ZN(g30290) );
NOR2_X4 U_g30291 ( .A1(g16460), .A2(g29987), .ZN(g30291) );
NOR2_X4 U_g30292 ( .A1(g13477), .A2(g29988), .ZN(g30292) );
NOR2_X4 U_g30293 ( .A1(g13480), .A2(g29989), .ZN(g30293) );
NOR2_X4 U_g30294 ( .A1(g13483), .A2(g29990), .ZN(g30294) );
NOR2_X4 U_g30295 ( .A1(g13485), .A2(g29991), .ZN(g30295) );
NOR2_X4 U_g30296 ( .A1(g13488), .A2(g29993), .ZN(g30296) );
NOR2_X4 U_g30297 ( .A1(g13490), .A2(g29994), .ZN(g30297) );
NOR2_X4 U_g30298 ( .A1(g13496), .A2(g29995), .ZN(g30298) );
NOR2_X4 U_g30299 ( .A1(g13499), .A2(g29996), .ZN(g30299) );
NOR2_X4 U_g30300 ( .A1(g13502), .A2(g30001), .ZN(g30300) );
NOR2_X4 U_g30301 ( .A1(g13504), .A2(g30002), .ZN(g30301) );
NOR2_X4 U_g30302 ( .A1(g13513), .A2(g30003), .ZN(g30302) );
NOR2_X4 U_g30303 ( .A1(g13516), .A2(g30005), .ZN(g30303) );
NOR2_X4 U_g30304 ( .A1(g13527), .A2(g30007), .ZN(g30304) );
NOR2_X4 U_g30338 ( .A1(g14297), .A2(g30225), .ZN(g30338) );
NOR2_X4 U_g30341 ( .A1(g14328), .A2(g30226), .ZN(g30341) );
NOR2_X4 U_g30356 ( .A1(g14419), .A2(g30227), .ZN(g30356) );
NOR2_X4 U_g30399 ( .A1(g30116), .A2(g30123), .ZN(g30399) );
NOR2_X4 U_g30400 ( .A1(g29997), .A2(g30127), .ZN(g30400) );
NOR2_X4 U_g30401 ( .A1(g29998), .A2(g30128), .ZN(g30401) );
NOR2_X4 U_g30402 ( .A1(g29999), .A2(g30129), .ZN(g30402) );
NOR2_X4 U_g30403 ( .A1(g30004), .A2(g30131), .ZN(g30403) );
NOR2_X4 U_g30404 ( .A1(g30006), .A2(g30132), .ZN(g30404) );
NOR2_X4 U_g30405 ( .A1(g30008), .A2(g30133), .ZN(g30405) );
NOR2_X4 U_g30406 ( .A1(g30009), .A2(g30138), .ZN(g30406) );
NOR2_X4 U_g30455 ( .A1(g13953), .A2(g30216), .ZN(g30455) );
NOR2_X4 U_g30468 ( .A1(g14007), .A2(g30217), .ZN(g30468) );
NOR2_X4 U_g30470 ( .A1(g14023), .A2(g30218), .ZN(g30470) );
NOR2_X4 U_g30482 ( .A1(g14067), .A2(g30219), .ZN(g30482) );
NOR2_X4 U_g30485 ( .A1(g14098), .A2(g30220), .ZN(g30485) );
NOR2_X4 U_g30487 ( .A1(g14114), .A2(g30221), .ZN(g30487) );
NOR2_X4 U_g30500 ( .A1(g14182), .A2(g30222), .ZN(g30500) );
NOR2_X4 U_g30503 ( .A1(g14213), .A2(g30223), .ZN(g30503) );
NOR2_X4 U_g30505 ( .A1(g14229), .A2(g30224), .ZN(g30505) );
NOR2_X4 U_g30566 ( .A1(g14327), .A2(g30398), .ZN(g30566) );
NOR2_X4 U_g30584 ( .A1(g30412), .A2(g2611), .ZN(g30584) );
NOR3_X4 U_g30588 ( .A1(g6119), .A2(g30412), .A3(g25353), .ZN(g30588) );
NOR2_X4 U_g30593 ( .A1(g30412), .A2(g2603), .ZN(g30593) );
NOR3_X4 U_g30594 ( .A1(g6119), .A2(g30412), .A3(g25419), .ZN(g30594) );
NOR3_X4 U_g30597 ( .A1(g6119), .A2(g30412), .A3(g25341), .ZN(g30597) );
NOR2_X4 U_g30601 ( .A1(g30412), .A2(g2604), .ZN(g30601) );
NOR3_X4 U_g30602 ( .A1(g6119), .A2(g30412), .A3(g25417), .ZN(g30602) );
NOR3_X4 U_g30605 ( .A1(g6119), .A2(g30412), .A3(g25333), .ZN(g30605) );
NOR2_X4 U_g30608 ( .A1(g30412), .A2(g2605), .ZN(g30608) );
NOR2_X4 U_g30609 ( .A1(g30412), .A2(g2606), .ZN(g30609) );
NOR3_X4 U_g30610 ( .A1(g6119), .A2(g30412), .A3(g25411), .ZN(g30610) );
NOR2_X4 U_g30613 ( .A1(g30412), .A2(g2607), .ZN(g30613) );
NOR3_X4 U_g30614 ( .A1(g6119), .A2(g30412), .A3(g25403), .ZN(g30614) );
NOR2_X4 U_g30617 ( .A1(g23850), .A2(g30412), .ZN(g30617) );
NOR2_X4 U_g30618 ( .A1(g30412), .A2(g25449), .ZN(g30618) );
NOR2_X4 U_g30621 ( .A1(g30412), .A2(g2608), .ZN(g30621) );
NOR3_X4 U_g30622 ( .A1(g6119), .A2(g30412), .A3(g25393), .ZN(g30622) );
NOR2_X4 U_g30625 ( .A1(g30412), .A2(g24660), .ZN(g30625) );
NOR2_X4 U_g30628 ( .A1(g30412), .A2(g2610), .ZN(g30628) );
NOR3_X4 U_g30629 ( .A1(g6119), .A2(g30412), .A3(g25378), .ZN(g30629) );
NOR3_X4 U_g30632 ( .A1(g6119), .A2(g30412), .A3(g25366), .ZN(g30632) );
NOR2_X4 U_g30635 ( .A1(g16108), .A2(g30407), .ZN(g30635) );
NOR2_X4 U_g30636 ( .A1(g16140), .A2(g30409), .ZN(g30636) );
NOR2_X4 U_g30637 ( .A1(g16141), .A2(g30410), .ZN(g30637) );
NOR2_X4 U_g30638 ( .A1(g16159), .A2(g30411), .ZN(g30638) );
NOR2_X4 U_g30639 ( .A1(g16186), .A2(g30436), .ZN(g30639) );
NOR2_X4 U_g30640 ( .A1(g16187), .A2(g30437), .ZN(g30640) );
NOR2_X4 U_g30641 ( .A1(g16188), .A2(g30438), .ZN(g30641) );
NOR2_X4 U_g30642 ( .A1(g16199), .A2(g30440), .ZN(g30642) );
NOR2_X4 U_g30643 ( .A1(g16200), .A2(g30441), .ZN(g30643) );
NOR2_X4 U_g30644 ( .A1(g16218), .A2(g30442), .ZN(g30644) );
NOR2_X4 U_g30645 ( .A1(g16240), .A2(g30444), .ZN(g30645) );
NOR2_X4 U_g30646 ( .A1(g16241), .A2(g30445), .ZN(g30646) );
NOR2_X4 U_g30647 ( .A1(g16251), .A2(g30447), .ZN(g30647) );
NOR2_X4 U_g30648 ( .A1(g16252), .A2(g30448), .ZN(g30648) );
NOR2_X4 U_g30649 ( .A1(g16253), .A2(g30449), .ZN(g30649) );
NOR2_X4 U_g30650 ( .A1(g16264), .A2(g30451), .ZN(g30650) );
NOR2_X4 U_g30651 ( .A1(g16265), .A2(g30452), .ZN(g30651) );
NOR2_X4 U_g30652 ( .A1(g16283), .A2(g30453), .ZN(g30652) );
NOR2_X4 U_g30653 ( .A1(g16289), .A2(g30454), .ZN(g30653) );
NOR2_X4 U_g30654 ( .A1(g16299), .A2(g30457), .ZN(g30654) );
NOR2_X4 U_g30655 ( .A1(g16300), .A2(g30458), .ZN(g30655) );
NOR2_X4 U_g30656 ( .A1(g16310), .A2(g30460), .ZN(g30656) );
NOR2_X4 U_g30657 ( .A1(g16311), .A2(g30461), .ZN(g30657) );
NOR2_X4 U_g30658 ( .A1(g16312), .A2(g30462), .ZN(g30658) );
NOR2_X4 U_g30659 ( .A1(g16323), .A2(g30464), .ZN(g30659) );
NOR2_X4 U_g30660 ( .A1(g16324), .A2(g30465), .ZN(g30660) );
NOR2_X4 U_g30661 ( .A1(g16345), .A2(g30467), .ZN(g30661) );
NOR2_X4 U_g30662 ( .A1(g16347), .A2(g30469), .ZN(g30662) );
NOR2_X4 U_g30663 ( .A1(g16357), .A2(g30472), .ZN(g30663) );
NOR2_X4 U_g30664 ( .A1(g16358), .A2(g30473), .ZN(g30664) );
NOR2_X4 U_g30665 ( .A1(g16368), .A2(g30475), .ZN(g30665) );
NOR2_X4 U_g30666 ( .A1(g16369), .A2(g30476), .ZN(g30666) );
NOR2_X4 U_g30667 ( .A1(g16370), .A2(g30477), .ZN(g30667) );
NOR2_X4 U_g30668 ( .A1(g16381), .A2(g30478), .ZN(g30668) );
NOR2_X4 U_g30669 ( .A1(g16383), .A2(g30481), .ZN(g30669) );
NOR2_X4 U_g30670 ( .A1(g16389), .A2(g30484), .ZN(g30670) );
NOR2_X4 U_g30671 ( .A1(g16391), .A2(g30486), .ZN(g30671) );
NOR2_X4 U_g30672 ( .A1(g16401), .A2(g30489), .ZN(g30672) );
NOR2_X4 U_g30673 ( .A1(g16402), .A2(g30490), .ZN(g30673) );
NOR2_X4 U_g30674 ( .A1(g16414), .A2(g30492), .ZN(g30674) );
NOR2_X4 U_g30675 ( .A1(g16416), .A2(g30495), .ZN(g30675) );
NOR2_X4 U_g30676 ( .A1(g16419), .A2(g30496), .ZN(g30676) );
NOR2_X4 U_g30677 ( .A1(g16421), .A2(g30499), .ZN(g30677) );
NOR2_X4 U_g30678 ( .A1(g16427), .A2(g30502), .ZN(g30678) );
NOR2_X4 U_g30679 ( .A1(g16429), .A2(g30504), .ZN(g30679) );
NOR2_X4 U_g30680 ( .A1(g16443), .A2(g30327), .ZN(g30680) );
NOR2_X4 U_g30681 ( .A1(g16448), .A2(g30330), .ZN(g30681) );
NOR2_X4 U_g30682 ( .A1(g16450), .A2(g30333), .ZN(g30682) );
NOR2_X4 U_g30683 ( .A1(g16453), .A2(g30334), .ZN(g30683) );
NOR2_X4 U_g30684 ( .A1(g16455), .A2(g30337), .ZN(g30684) );
NOR3_X4 U_g30685 ( .A1(g29992), .A2(g30000), .A3(g30372), .ZN(g30685) );
NOR2_X4 U_g30686 ( .A1(g16461), .A2(g30340), .ZN(g30686) );
NOR2_X4 U_g30687 ( .A1(g13479), .A2(g30345), .ZN(g30687) );
NOR2_X4 U_g30688 ( .A1(g13484), .A2(g30348), .ZN(g30688) );
NOR2_X4 U_g30689 ( .A1(g13486), .A2(g30351), .ZN(g30689) );
NOR2_X4 U_g30690 ( .A1(g13489), .A2(g30352), .ZN(g30690) );
NOR2_X4 U_g30691 ( .A1(g13491), .A2(g30355), .ZN(g30691) );
NOR2_X4 U_g30692 ( .A1(g13498), .A2(g30361), .ZN(g30692) );
NOR2_X4 U_g30693 ( .A1(g13503), .A2(g30364), .ZN(g30693) );
NOR2_X4 U_g30694 ( .A1(g13505), .A2(g30367), .ZN(g30694) );
NOR2_X4 U_g30695 ( .A1(g13515), .A2(g30374), .ZN(g30695) );
NOR2_X4 U_g30699 ( .A1(g13914), .A2(g30387), .ZN(g30699) );
NOR2_X4 U_g30700 ( .A1(g13952), .A2(g30388), .ZN(g30700) );
NOR2_X4 U_g30701 ( .A1(g13970), .A2(g30389), .ZN(g30701) );
NOR2_X4 U_g30702 ( .A1(g14006), .A2(g30390), .ZN(g30702) );
NOR2_X4 U_g30703 ( .A1(g14022), .A2(g30391), .ZN(g30703) );
NOR2_X4 U_g30704 ( .A1(g14040), .A2(g30392), .ZN(g30704) );
NOR2_X4 U_g30705 ( .A1(g14097), .A2(g30393), .ZN(g30705) );
NOR2_X4 U_g30706 ( .A1(g14113), .A2(g30394), .ZN(g30706) );
NOR2_X4 U_g30707 ( .A1(g14131), .A2(g30395), .ZN(g30707) );
NOR2_X4 U_g30708 ( .A1(g14212), .A2(g30396), .ZN(g30708) );
NOR2_X4 U_g30709 ( .A1(g14228), .A2(g30397), .ZN(g30709) );
NOR2_X4 U_g30780 ( .A1(g30625), .A2(g22387), .ZN(g30780) );
NOR2_X4 U_g30783 ( .A1(g30618), .A2(g22387), .ZN(g30783) );
NOR2_X4 U_g30785 ( .A1(g30618), .A2(g22387), .ZN(g30785) );
NOR2_X4 U_g30786 ( .A1(g30625), .A2(g22387), .ZN(g30786) );
NOR2_X4 U_g30787 ( .A1(g30594), .A2(g22387), .ZN(g30787) );
NOR2_X4 U_g30788 ( .A1(g30602), .A2(g22387), .ZN(g30788) );
NOR2_X4 U_g30789 ( .A1(g30575), .A2(g22387), .ZN(g30789) );
NOR2_X4 U_g30790 ( .A1(g30575), .A2(g22387), .ZN(g30790) );
NOR2_X4 U_g30796 ( .A1(g16069), .A2(g30696), .ZN(g30796) );
NOR2_X4 U_g30798 ( .A1(g16134), .A2(g30697), .ZN(g30798) );
NOR2_X4 U_g30801 ( .A1(g16237), .A2(g30698), .ZN(g30801) );
NOR2_X4 U_g30929 ( .A1(g30728), .A2(g30736), .ZN(g30929) );
NOR2_X4 U_g30930 ( .A1(g30735), .A2(g30744), .ZN(g30930) );
NOR2_X4 U_g30931 ( .A1(g30743), .A2(g30750), .ZN(g30931) );
NOR2_X4 U_g30932 ( .A1(g30754), .A2(g30757), .ZN(g30932) );
NOR2_X4 U_g30933 ( .A1(g30755), .A2(g30758), .ZN(g30933) );
NOR2_X4 U_g30934 ( .A1(g30759), .A2(g30761), .ZN(g30934) );
NOR2_X4 U_g30935 ( .A1(g30760), .A2(g30762), .ZN(g30935) );
NOR2_X4 U_g30936 ( .A1(g30763), .A2(g30764), .ZN(g30936) );
NOR2_X4 U_g30954 ( .A1(g30916), .A2(g30944), .ZN(g30954) );
NOR2_X4 U_g30955 ( .A1(g30918), .A2(g30945), .ZN(g30955) );
NOR2_X4 U_g30956 ( .A1(g30919), .A2(g30946), .ZN(g30956) );
NOR2_X4 U_g30957 ( .A1(g30920), .A2(g30947), .ZN(g30957) );
NOR2_X4 U_g30958 ( .A1(g30922), .A2(g30948), .ZN(g30958) );
NOR2_X4 U_g30959 ( .A1(g30923), .A2(g30949), .ZN(g30959) );
NOR2_X4 U_g30960 ( .A1(g30924), .A2(g30950), .ZN(g30960) );
NOR2_X4 U_g30961 ( .A1(g30925), .A2(g30951), .ZN(g30961) );
NOR3_X4 U_g30970 ( .A1(g30917), .A2(g30921), .A3(g30953), .ZN(g30970) );

DFF_X2 U_g2814 ( .D(g16475), .Q(g2814), .CK(CK) );
DFF_X2 U_g2817 ( .D(g20571), .Q(g2817), .CK(CK) );
DFF_X2 U_g2933 ( .D(g20588), .Q(g2933), .CK(CK) );
DFF_X2 U_g2950 ( .D(g21951), .Q(g2950), .CK(CK) );
DFF_X2 U_g2883 ( .D(g23315), .Q(g2883), .CK(CK) );
DFF_X2 U_g2888 ( .D(g24423), .Q(g2888), .CK(CK) );
DFF_X2 U_g2896 ( .D(g25175), .Q(g2896), .CK(CK) );
DFF_X2 U_g2892 ( .D(g26019), .Q(g2892), .CK(CK) );
DFF_X2 U_g2903 ( .D(g26747), .Q(g2903), .CK(CK) );
DFF_X2 U_g2900 ( .D(g27237), .Q(g2900), .CK(CK) );
DFF_X2 U_g2908 ( .D(g27715), .Q(g2908), .CK(CK) );
DFF_X2 U_g2912 ( .D(g24424), .Q(g2912), .CK(CK) );
DFF_X2 U_g2917 ( .D(g25174), .Q(g2917), .CK(CK) );
DFF_X2 U_g2924 ( .D(g26020), .Q(g2924), .CK(CK) );
DFF_X2 U_g2920 ( .D(g26746), .Q(g2920), .CK(CK) );
DFF_X2 U_g2984 ( .D(g19061), .Q(g2984), .CK(CK) );
DFF_X2 U_g2985 ( .D(g19060), .Q(g2985), .CK(CK) );
DFF_X2 U_g2930 ( .D(g19062), .Q(g2930), .CK(CK) );
DFF_X2 U_g2929 ( .D(g2930), .Q(g2929), .CK(CK) );
DFF_X2 U_g2879 ( .D(g16494), .Q(g2879), .CK(CK) );
DFF_X2 U_g2934 ( .D(g16476), .Q(g2934), .CK(CK) );
DFF_X2 U_g2935 ( .D(g16477), .Q(g2935), .CK(CK) );
DFF_X2 U_g2938 ( .D(g16478), .Q(g2938), .CK(CK) );
DFF_X2 U_g2941 ( .D(g16479), .Q(g2941), .CK(CK) );
DFF_X2 U_g2944 ( .D(g16480), .Q(g2944), .CK(CK) );
DFF_X2 U_g2947 ( .D(g16481), .Q(g2947), .CK(CK) );
DFF_X2 U_g2953 ( .D(g16482), .Q(g2953), .CK(CK) );
DFF_X2 U_g2956 ( .D(g16483), .Q(g2956), .CK(CK) );
DFF_X2 U_g2959 ( .D(g16484), .Q(g2959), .CK(CK) );
DFF_X2 U_g2962 ( .D(g16485), .Q(g2962), .CK(CK) );
DFF_X2 U_g2963 ( .D(g16486), .Q(g2963), .CK(CK) );
DFF_X2 U_g2966 ( .D(g16487), .Q(g2966), .CK(CK) );
DFF_X2 U_g2969 ( .D(g16488), .Q(g2969), .CK(CK) );
DFF_X2 U_g2972 ( .D(g16489), .Q(g2972), .CK(CK) );
DFF_X2 U_g2975 ( .D(g16490), .Q(g2975), .CK(CK) );
DFF_X2 U_g2978 ( .D(g16491), .Q(g2978), .CK(CK) );
DFF_X2 U_g2981 ( .D(g16492), .Q(g2981), .CK(CK) );
DFF_X2 U_g2874 ( .D(g16493), .Q(g2874), .CK(CK) );
DFF_X2 U_g1506 ( .D(g20572), .Q(g1506), .CK(CK) );
DFF_X2 U_g1501 ( .D(g20573), .Q(g1501), .CK(CK) );
DFF_X2 U_g1496 ( .D(g20574), .Q(g1496), .CK(CK) );
DFF_X2 U_g1491 ( .D(g20575), .Q(g1491), .CK(CK) );
DFF_X2 U_g1486 ( .D(g20576), .Q(g1486), .CK(CK) );
DFF_X2 U_g1481 ( .D(g20577), .Q(g1481), .CK(CK) );
DFF_X2 U_g1476 ( .D(g20578), .Q(g1476), .CK(CK) );
DFF_X2 U_g1471 ( .D(g20579), .Q(g1471), .CK(CK) );
DFF_X2 U_g2877 ( .D(g23313), .Q(g2877), .CK(CK) );
DFF_X2 U_g2861 ( .D(g21960), .Q(g2861), .CK(CK) );
DFF_X2 U_g813 ( .D(g2861), .Q(g813), .CK(CK) );
DFF_X2 U_g2864 ( .D(g21961), .Q(g2864), .CK(CK) );
DFF_X2 U_g809 ( .D(g2864), .Q(g809), .CK(CK) );
DFF_X2 U_g2867 ( .D(g21962), .Q(g2867), .CK(CK) );
DFF_X2 U_g805 ( .D(g2867), .Q(g805), .CK(CK) );
DFF_X2 U_g2870 ( .D(g21963), .Q(g2870), .CK(CK) );
DFF_X2 U_g801 ( .D(g2870), .Q(g801), .CK(CK) );
DFF_X2 U_g2818 ( .D(g21947), .Q(g2818), .CK(CK) );
DFF_X2 U_g797 ( .D(g2818), .Q(g797), .CK(CK) );
DFF_X2 U_g2821 ( .D(g21948), .Q(g2821), .CK(CK) );
DFF_X2 U_g793 ( .D(g2821), .Q(g793), .CK(CK) );
DFF_X2 U_g2824 ( .D(g21949), .Q(g2824), .CK(CK) );
DFF_X2 U_g789 ( .D(g2824), .Q(g789), .CK(CK) );
DFF_X2 U_g2827 ( .D(g21950), .Q(g2827), .CK(CK) );
DFF_X2 U_g785 ( .D(g2827), .Q(g785), .CK(CK) );
DFF_X2 U_g2830 ( .D(g23312), .Q(g2830), .CK(CK) );
DFF_X2 U_g2873 ( .D(g2830), .Q(g2873), .CK(CK) );
DFF_X2 U_g2833 ( .D(g21952), .Q(g2833), .CK(CK) );
DFF_X2 U_g125 ( .D(g2833), .Q(g125), .CK(CK) );
DFF_X2 U_g2836 ( .D(g21953), .Q(g2836), .CK(CK) );
DFF_X2 U_g121 ( .D(g2836), .Q(g121), .CK(CK) );
DFF_X2 U_g2839 ( .D(g21954), .Q(g2839), .CK(CK) );
DFF_X2 U_g117 ( .D(g2839), .Q(g117), .CK(CK) );
DFF_X2 U_g2842 ( .D(g21955), .Q(g2842), .CK(CK) );
DFF_X2 U_g113 ( .D(g2842), .Q(g113), .CK(CK) );
DFF_X2 U_g2845 ( .D(g21956), .Q(g2845), .CK(CK) );
DFF_X2 U_g109 ( .D(g2845), .Q(g109), .CK(CK) );
DFF_X2 U_g2848 ( .D(g21957), .Q(g2848), .CK(CK) );
DFF_X2 U_g105 ( .D(g2848), .Q(g105), .CK(CK) );
DFF_X2 U_g2851 ( .D(g21958), .Q(g2851), .CK(CK) );
DFF_X2 U_g101 ( .D(g2851), .Q(g101), .CK(CK) );
DFF_X2 U_g2854 ( .D(g21959), .Q(g2854), .CK(CK) );
DFF_X2 U_g97 ( .D(g2854), .Q(g97), .CK(CK) );
DFF_X2 U_g2858 ( .D(g23316), .Q(g2858), .CK(CK) );
DFF_X2 U_g2857 ( .D(g2858), .Q(g2857), .CK(CK) );
DFF_X2 U_g2200 ( .D(g20587), .Q(g2200), .CK(CK) );
DFF_X2 U_g2195 ( .D(g20585), .Q(g2195), .CK(CK) );
DFF_X2 U_g2190 ( .D(g20586), .Q(g2190), .CK(CK) );
DFF_X2 U_g2185 ( .D(g20584), .Q(g2185), .CK(CK) );
DFF_X2 U_g2180 ( .D(g20583), .Q(g2180), .CK(CK) );
DFF_X2 U_g2175 ( .D(g20582), .Q(g2175), .CK(CK) );
DFF_X2 U_g2170 ( .D(g20581), .Q(g2170), .CK(CK) );
DFF_X2 U_g2165 ( .D(g20580), .Q(g2165), .CK(CK) );
DFF_X2 U_g2878 ( .D(g23314), .Q(g2878), .CK(CK) );
DFF_X2 U_g3129 ( .D(g13475), .Q(g3129), .CK(CK) );
DFF_X2 U_g3117 ( .D(g3129), .Q(g3117), .CK(CK) );
DFF_X2 U_g3109 ( .D(g3117), .Q(g3109), .CK(CK) );
DFF_X2 U_g3210 ( .D(g20630), .Q(g3210), .CK(CK) );
DFF_X2 U_g3211 ( .D(g20631), .Q(g3211), .CK(CK) );
DFF_X2 U_g3084 ( .D(g20632), .Q(g3084), .CK(CK) );
DFF_X2 U_g3085 ( .D(g20609), .Q(g3085), .CK(CK) );
DFF_X2 U_g3086 ( .D(g20610), .Q(g3086), .CK(CK) );
DFF_X2 U_g3087 ( .D(g20611), .Q(g3087), .CK(CK) );
DFF_X2 U_g3091 ( .D(g20612), .Q(g3091), .CK(CK) );
DFF_X2 U_g3092 ( .D(g20613), .Q(g3092), .CK(CK) );
DFF_X2 U_g3093 ( .D(g20614), .Q(g3093), .CK(CK) );
DFF_X2 U_g3094 ( .D(g20615), .Q(g3094), .CK(CK) );
DFF_X2 U_g3095 ( .D(g20616), .Q(g3095), .CK(CK) );
DFF_X2 U_g3096 ( .D(g20617), .Q(g3096), .CK(CK) );
DFF_X2 U_g3097 ( .D(g26751), .Q(g3097), .CK(CK) );
DFF_X2 U_g3098 ( .D(g26752), .Q(g3098), .CK(CK) );
DFF_X2 U_g3099 ( .D(g26753), .Q(g3099), .CK(CK) );
DFF_X2 U_g3100 ( .D(g29163), .Q(g3100), .CK(CK) );
DFF_X2 U_g3101 ( .D(g29164), .Q(g3101), .CK(CK) );
DFF_X2 U_g3102 ( .D(g29165), .Q(g3102), .CK(CK) );
DFF_X2 U_g3103 ( .D(g30120), .Q(g3103), .CK(CK) );
DFF_X2 U_g3104 ( .D(g30121), .Q(g3104), .CK(CK) );
DFF_X2 U_g3105 ( .D(g30122), .Q(g3105), .CK(CK) );
DFF_X2 U_g3106 ( .D(g30941), .Q(g3106), .CK(CK) );
DFF_X2 U_g3107 ( .D(g30942), .Q(g3107), .CK(CK) );
DFF_X2 U_g3108 ( .D(g30943), .Q(g3108), .CK(CK) );
DFF_X2 U_g3155 ( .D(g20618), .Q(g3155), .CK(CK) );
DFF_X2 U_g3158 ( .D(g20619), .Q(g3158), .CK(CK) );
DFF_X2 U_g3161 ( .D(g20620), .Q(g3161), .CK(CK) );
DFF_X2 U_g3164 ( .D(g20621), .Q(g3164), .CK(CK) );
DFF_X2 U_g3167 ( .D(g20622), .Q(g3167), .CK(CK) );
DFF_X2 U_g3170 ( .D(g20623), .Q(g3170), .CK(CK) );
DFF_X2 U_g3173 ( .D(g20624), .Q(g3173), .CK(CK) );
DFF_X2 U_g3176 ( .D(g20625), .Q(g3176), .CK(CK) );
DFF_X2 U_g3179 ( .D(g20626), .Q(g3179), .CK(CK) );
DFF_X2 U_g3182 ( .D(g20627), .Q(g3182), .CK(CK) );
DFF_X2 U_g3185 ( .D(g20628), .Q(g3185), .CK(CK) );
DFF_X2 U_g3088 ( .D(g20629), .Q(g3088), .CK(CK) );
DFF_X2 U_g3191 ( .D(g27717), .Q(g3191), .CK(CK) );
DFF_X2 U_g3194 ( .D(g28316), .Q(g3194), .CK(CK) );
DFF_X2 U_g3197 ( .D(g28317), .Q(g3197), .CK(CK) );
DFF_X2 U_g3198 ( .D(g28318), .Q(g3198), .CK(CK) );
DFF_X2 U_g3201 ( .D(g28704), .Q(g3201), .CK(CK) );
DFF_X2 U_g3204 ( .D(g28705), .Q(g3204), .CK(CK) );
DFF_X2 U_g3207 ( .D(g28706), .Q(g3207), .CK(CK) );
DFF_X2 U_g3188 ( .D(g29463), .Q(g3188), .CK(CK) );
DFF_X2 U_g3133 ( .D(g29656), .Q(g3133), .CK(CK) );
DFF_X2 U_g3132 ( .D(g28698), .Q(g3132), .CK(CK) );
DFF_X2 U_g3128 ( .D(g29166), .Q(g3128), .CK(CK) );
DFF_X2 U_g3127 ( .D(g28697), .Q(g3127), .CK(CK) );
DFF_X2 U_g3126 ( .D(g28315), .Q(g3126), .CK(CK) );
DFF_X2 U_g3125 ( .D(g28696), .Q(g3125), .CK(CK) );
DFF_X2 U_g3124 ( .D(g28314), .Q(g3124), .CK(CK) );
DFF_X2 U_g3123 ( .D(g28313), .Q(g3123), .CK(CK) );
DFF_X2 U_g3120 ( .D(g28695), .Q(g3120), .CK(CK) );
DFF_X2 U_g3114 ( .D(g28694), .Q(g3114), .CK(CK) );
DFF_X2 U_g3113 ( .D(g28693), .Q(g3113), .CK(CK) );
DFF_X2 U_g3112 ( .D(g28312), .Q(g3112), .CK(CK) );
DFF_X2 U_g3110 ( .D(g28311), .Q(g3110), .CK(CK) );
DFF_X2 U_g3111 ( .D(g28310), .Q(g3111), .CK(CK) );
DFF_X2 U_g3139 ( .D(g29461), .Q(g3139), .CK(CK) );
DFF_X2 U_g3136 ( .D(g28701), .Q(g3136), .CK(CK) );
DFF_X2 U_g3134 ( .D(g28700), .Q(g3134), .CK(CK) );
DFF_X2 U_g3135 ( .D(g28699), .Q(g3135), .CK(CK) );
DFF_X2 U_g3151 ( .D(g29462), .Q(g3151), .CK(CK) );
DFF_X2 U_g3142 ( .D(g28703), .Q(g3142), .CK(CK) );
DFF_X2 U_g3147 ( .D(g28702), .Q(g3147), .CK(CK) );
DFF_X2 U_g185 ( .D(g29657), .Q(g185), .CK(CK) );
DFF_X2 U_g138 ( .D(g13405), .Q(g138), .CK(CK) );
DFF_X2 U_g135 ( .D(g138), .Q(g135), .CK(CK) );
DFF_X2 U_g165 ( .D(g135), .Q(g165), .CK(CK) );
DFF_X2 U_g130 ( .D(g24259), .Q(g130), .CK(CK) );
DFF_X2 U_g131 ( .D(g24260), .Q(g131), .CK(CK) );
DFF_X2 U_g129 ( .D(g24261), .Q(g129), .CK(CK) );
DFF_X2 U_g133 ( .D(g24262), .Q(g133), .CK(CK) );
DFF_X2 U_g134 ( .D(g24263), .Q(g134), .CK(CK) );
DFF_X2 U_g132 ( .D(g24264), .Q(g132), .CK(CK) );
DFF_X2 U_g142 ( .D(g24265), .Q(g142), .CK(CK) );
DFF_X2 U_g143 ( .D(g24266), .Q(g143), .CK(CK) );
DFF_X2 U_g141 ( .D(g24267), .Q(g141), .CK(CK) );
DFF_X2 U_g145 ( .D(g24268), .Q(g145), .CK(CK) );
DFF_X2 U_g146 ( .D(g24269), .Q(g146), .CK(CK) );
DFF_X2 U_g144 ( .D(g24270), .Q(g144), .CK(CK) );
DFF_X2 U_g148 ( .D(g24271), .Q(g148), .CK(CK) );
DFF_X2 U_g149 ( .D(g24272), .Q(g149), .CK(CK) );
DFF_X2 U_g147 ( .D(g24273), .Q(g147), .CK(CK) );
DFF_X2 U_g151 ( .D(g24274), .Q(g151), .CK(CK) );
DFF_X2 U_g152 ( .D(g24275), .Q(g152), .CK(CK) );
DFF_X2 U_g150 ( .D(g24276), .Q(g150), .CK(CK) );
DFF_X2 U_g154 ( .D(g24277), .Q(g154), .CK(CK) );
DFF_X2 U_g155 ( .D(g24278), .Q(g155), .CK(CK) );
DFF_X2 U_g153 ( .D(g24279), .Q(g153), .CK(CK) );
DFF_X2 U_g157 ( .D(g24280), .Q(g157), .CK(CK) );
DFF_X2 U_g158 ( .D(g24281), .Q(g158), .CK(CK) );
DFF_X2 U_g156 ( .D(g24282), .Q(g156), .CK(CK) );
DFF_X2 U_g160 ( .D(g24283), .Q(g160), .CK(CK) );
DFF_X2 U_g161 ( .D(g24284), .Q(g161), .CK(CK) );
DFF_X2 U_g159 ( .D(g24285), .Q(g159), .CK(CK) );
DFF_X2 U_g163 ( .D(g24286), .Q(g163), .CK(CK) );
DFF_X2 U_g164 ( .D(g24287), .Q(g164), .CK(CK) );
DFF_X2 U_g162 ( .D(g24288), .Q(g162), .CK(CK) );
DFF_X2 U_g169 ( .D(g26679), .Q(g169), .CK(CK) );
DFF_X2 U_g170 ( .D(g26680), .Q(g170), .CK(CK) );
DFF_X2 U_g168 ( .D(g26681), .Q(g168), .CK(CK) );
DFF_X2 U_g172 ( .D(g26682), .Q(g172), .CK(CK) );
DFF_X2 U_g173 ( .D(g26683), .Q(g173), .CK(CK) );
DFF_X2 U_g171 ( .D(g26684), .Q(g171), .CK(CK) );
DFF_X2 U_g175 ( .D(g26685), .Q(g175), .CK(CK) );
DFF_X2 U_g176 ( .D(g26686), .Q(g176), .CK(CK) );
DFF_X2 U_g174 ( .D(g26687), .Q(g174), .CK(CK) );
DFF_X2 U_g178 ( .D(g26688), .Q(g178), .CK(CK) );
DFF_X2 U_g179 ( .D(g26689), .Q(g179), .CK(CK) );
DFF_X2 U_g177 ( .D(g26690), .Q(g177), .CK(CK) );
DFF_X2 U_g186 ( .D(g30506), .Q(g186), .CK(CK) );
DFF_X2 U_g189 ( .D(g30507), .Q(g189), .CK(CK) );
DFF_X2 U_g192 ( .D(g30508), .Q(g192), .CK(CK) );
DFF_X2 U_g231 ( .D(g30842), .Q(g231), .CK(CK) );
DFF_X2 U_g234 ( .D(g30843), .Q(g234), .CK(CK) );
DFF_X2 U_g237 ( .D(g30844), .Q(g237), .CK(CK) );
DFF_X2 U_g195 ( .D(g30836), .Q(g195), .CK(CK) );
DFF_X2 U_g198 ( .D(g30837), .Q(g198), .CK(CK) );
DFF_X2 U_g201 ( .D(g30838), .Q(g201), .CK(CK) );
DFF_X2 U_g240 ( .D(g30845), .Q(g240), .CK(CK) );
DFF_X2 U_g243 ( .D(g30846), .Q(g243), .CK(CK) );
DFF_X2 U_g246 ( .D(g30847), .Q(g246), .CK(CK) );
DFF_X2 U_g204 ( .D(g30509), .Q(g204), .CK(CK) );
DFF_X2 U_g207 ( .D(g30510), .Q(g207), .CK(CK) );
DFF_X2 U_g210 ( .D(g30511), .Q(g210), .CK(CK) );
DFF_X2 U_g249 ( .D(g30515), .Q(g249), .CK(CK) );
DFF_X2 U_g252 ( .D(g30516), .Q(g252), .CK(CK) );
DFF_X2 U_g255 ( .D(g30517), .Q(g255), .CK(CK) );
DFF_X2 U_g213 ( .D(g30512), .Q(g213), .CK(CK) );
DFF_X2 U_g216 ( .D(g30513), .Q(g216), .CK(CK) );
DFF_X2 U_g219 ( .D(g30514), .Q(g219), .CK(CK) );
DFF_X2 U_g258 ( .D(g30518), .Q(g258), .CK(CK) );
DFF_X2 U_g261 ( .D(g30519), .Q(g261), .CK(CK) );
DFF_X2 U_g264 ( .D(g30520), .Q(g264), .CK(CK) );
DFF_X2 U_g222 ( .D(g30839), .Q(g222), .CK(CK) );
DFF_X2 U_g225 ( .D(g30840), .Q(g225), .CK(CK) );
DFF_X2 U_g228 ( .D(g30841), .Q(g228), .CK(CK) );
DFF_X2 U_g267 ( .D(g30848), .Q(g267), .CK(CK) );
DFF_X2 U_g270 ( .D(g30849), .Q(g270), .CK(CK) );
DFF_X2 U_g273 ( .D(g30850), .Q(g273), .CK(CK) );
DFF_X2 U_g92 ( .D(g25983), .Q(g92), .CK(CK) );
DFF_X2 U_g88 ( .D(g26678), .Q(g88), .CK(CK) );
DFF_X2 U_g83 ( .D(g27189), .Q(g83), .CK(CK) );
DFF_X2 U_g79 ( .D(g27683), .Q(g79), .CK(CK) );
DFF_X2 U_g74 ( .D(g28206), .Q(g74), .CK(CK) );
DFF_X2 U_g70 ( .D(g28673), .Q(g70), .CK(CK) );
DFF_X2 U_g65 ( .D(g29131), .Q(g65), .CK(CK) );
DFF_X2 U_g61 ( .D(g29413), .Q(g61), .CK(CK) );
DFF_X2 U_g56 ( .D(g29627), .Q(g56), .CK(CK) );
DFF_X2 U_g52 ( .D(g29794), .Q(g52), .CK(CK) );
DFF_X2 U_g180 ( .D(g20555), .Q(g180), .CK(CK) );
DFF_X2 U_g182 ( .D(g180), .Q(g182), .CK(CK) );
DFF_X2 U_g181 ( .D(g182), .Q(g181), .CK(CK) );
DFF_X2 U_g276 ( .D(g13406), .Q(g276), .CK(CK) );
DFF_X2 U_g405 ( .D(g276), .Q(g405), .CK(CK) );
DFF_X2 U_g401 ( .D(g405), .Q(g401), .CK(CK) );
DFF_X2 U_g309 ( .D(g11496), .Q(g309), .CK(CK) );
DFF_X2 U_g354 ( .D(g28207), .Q(g354), .CK(CK) );
DFF_X2 U_g343 ( .D(g28208), .Q(g343), .CK(CK) );
DFF_X2 U_g346 ( .D(g28209), .Q(g346), .CK(CK) );
DFF_X2 U_g369 ( .D(g28210), .Q(g369), .CK(CK) );
DFF_X2 U_g358 ( .D(g28211), .Q(g358), .CK(CK) );
DFF_X2 U_g361 ( .D(g28212), .Q(g361), .CK(CK) );
DFF_X2 U_g384 ( .D(g28213), .Q(g384), .CK(CK) );
DFF_X2 U_g373 ( .D(g28214), .Q(g373), .CK(CK) );
DFF_X2 U_g376 ( .D(g28215), .Q(g376), .CK(CK) );
DFF_X2 U_g398 ( .D(g28216), .Q(g398), .CK(CK) );
DFF_X2 U_g388 ( .D(g28217), .Q(g388), .CK(CK) );
DFF_X2 U_g391 ( .D(g28218), .Q(g391), .CK(CK) );
DFF_X2 U_g408 ( .D(g29414), .Q(g408), .CK(CK) );
DFF_X2 U_g411 ( .D(g29415), .Q(g411), .CK(CK) );
DFF_X2 U_g414 ( .D(g29416), .Q(g414), .CK(CK) );
DFF_X2 U_g417 ( .D(g29631), .Q(g417), .CK(CK) );
DFF_X2 U_g420 ( .D(g29632), .Q(g420), .CK(CK) );
DFF_X2 U_g423 ( .D(g29633), .Q(g423), .CK(CK) );
DFF_X2 U_g427 ( .D(g29417), .Q(g427), .CK(CK) );
DFF_X2 U_g428 ( .D(g29418), .Q(g428), .CK(CK) );
DFF_X2 U_g426 ( .D(g29419), .Q(g426), .CK(CK) );
DFF_X2 U_g429 ( .D(g27684), .Q(g429), .CK(CK) );
DFF_X2 U_g432 ( .D(g27685), .Q(g432), .CK(CK) );
DFF_X2 U_g435 ( .D(g27686), .Q(g435), .CK(CK) );
DFF_X2 U_g438 ( .D(g27687), .Q(g438), .CK(CK) );
DFF_X2 U_g441 ( .D(g27688), .Q(g441), .CK(CK) );
DFF_X2 U_g444 ( .D(g27689), .Q(g444), .CK(CK) );
DFF_X2 U_g448 ( .D(g28674), .Q(g448), .CK(CK) );
DFF_X2 U_g449 ( .D(g28675), .Q(g449), .CK(CK) );
DFF_X2 U_g447 ( .D(g28676), .Q(g447), .CK(CK) );
DFF_X2 U_g312 ( .D(g29795), .Q(g312), .CK(CK) );
DFF_X2 U_g313 ( .D(g29796), .Q(g313), .CK(CK) );
DFF_X2 U_g314 ( .D(g29797), .Q(g314), .CK(CK) );
DFF_X2 U_g315 ( .D(g30851), .Q(g315), .CK(CK) );
DFF_X2 U_g316 ( .D(g30852), .Q(g316), .CK(CK) );
DFF_X2 U_g317 ( .D(g30853), .Q(g317), .CK(CK) );
DFF_X2 U_g318 ( .D(g30710), .Q(g318), .CK(CK) );
DFF_X2 U_g319 ( .D(g30711), .Q(g319), .CK(CK) );
DFF_X2 U_g320 ( .D(g30712), .Q(g320), .CK(CK) );
DFF_X2 U_g322 ( .D(g29628), .Q(g322), .CK(CK) );
DFF_X2 U_g323 ( .D(g29629), .Q(g323), .CK(CK) );
DFF_X2 U_g321 ( .D(g29630), .Q(g321), .CK(CK) );
DFF_X2 U_g403 ( .D(g27191), .Q(g403), .CK(CK) );
DFF_X2 U_g404 ( .D(g27192), .Q(g404), .CK(CK) );
DFF_X2 U_g402 ( .D(g27193), .Q(g402), .CK(CK) );
DFF_X2 U_g450 ( .D(g11509), .Q(g450), .CK(CK) );
DFF_X2 U_g451 ( .D(g450), .Q(g451), .CK(CK) );
DFF_X2 U_g452 ( .D(g11510), .Q(g452), .CK(CK) );
DFF_X2 U_g453 ( .D(g452), .Q(g453), .CK(CK) );
DFF_X2 U_g454 ( .D(g11511), .Q(g454), .CK(CK) );
DFF_X2 U_g279 ( .D(g454), .Q(g279), .CK(CK) );
DFF_X2 U_g280 ( .D(g11491), .Q(g280), .CK(CK) );
DFF_X2 U_g281 ( .D(g280), .Q(g281), .CK(CK) );
DFF_X2 U_g282 ( .D(g11492), .Q(g282), .CK(CK) );
DFF_X2 U_g283 ( .D(g282), .Q(g283), .CK(CK) );
DFF_X2 U_g284 ( .D(g11493), .Q(g284), .CK(CK) );
DFF_X2 U_g285 ( .D(g284), .Q(g285), .CK(CK) );
DFF_X2 U_g286 ( .D(g11494), .Q(g286), .CK(CK) );
DFF_X2 U_g287 ( .D(g286), .Q(g287), .CK(CK) );
DFF_X2 U_g288 ( .D(g11495), .Q(g288), .CK(CK) );
DFF_X2 U_g289 ( .D(g288), .Q(g289), .CK(CK) );
DFF_X2 U_g290 ( .D(g13407), .Q(g290), .CK(CK) );
DFF_X2 U_g291 ( .D(g290), .Q(g291), .CK(CK) );
DFF_X2 U_g299 ( .D(g19012), .Q(g299), .CK(CK) );
DFF_X2 U_g305 ( .D(g23148), .Q(g305), .CK(CK) );
DFF_X2 U_g308 ( .D(g23149), .Q(g308), .CK(CK) );
DFF_X2 U_g297 ( .D(g23150), .Q(g297), .CK(CK) );
DFF_X2 U_g296 ( .D(g23151), .Q(g296), .CK(CK) );
DFF_X2 U_g295 ( .D(g23152), .Q(g295), .CK(CK) );
DFF_X2 U_g294 ( .D(g23153), .Q(g294), .CK(CK) );
DFF_X2 U_g304 ( .D(g19016), .Q(g304), .CK(CK) );
DFF_X2 U_g303 ( .D(g19015), .Q(g303), .CK(CK) );
DFF_X2 U_g302 ( .D(g19014), .Q(g302), .CK(CK) );
DFF_X2 U_g301 ( .D(g19013), .Q(g301), .CK(CK) );
DFF_X2 U_g300 ( .D(g25130), .Q(g300), .CK(CK) );
DFF_X2 U_g298 ( .D(g27190), .Q(g298), .CK(CK) );
DFF_X2 U_g342 ( .D(g11497), .Q(g342), .CK(CK) );
DFF_X2 U_g349 ( .D(g342), .Q(g349), .CK(CK) );
DFF_X2 U_g350 ( .D(g11498), .Q(g350), .CK(CK) );
DFF_X2 U_g351 ( .D(g350), .Q(g351), .CK(CK) );
DFF_X2 U_g352 ( .D(g11499), .Q(g352), .CK(CK) );
DFF_X2 U_g353 ( .D(g352), .Q(g353), .CK(CK) );
DFF_X2 U_g357 ( .D(g11500), .Q(g357), .CK(CK) );
DFF_X2 U_g364 ( .D(g357), .Q(g364), .CK(CK) );
DFF_X2 U_g365 ( .D(g11501), .Q(g365), .CK(CK) );
DFF_X2 U_g366 ( .D(g365), .Q(g366), .CK(CK) );
DFF_X2 U_g367 ( .D(g11502), .Q(g367), .CK(CK) );
DFF_X2 U_g368 ( .D(g367), .Q(g368), .CK(CK) );
DFF_X2 U_g372 ( .D(g11503), .Q(g372), .CK(CK) );
DFF_X2 U_g379 ( .D(g372), .Q(g379), .CK(CK) );
DFF_X2 U_g380 ( .D(g11504), .Q(g380), .CK(CK) );
DFF_X2 U_g381 ( .D(g380), .Q(g381), .CK(CK) );
DFF_X2 U_g382 ( .D(g11505), .Q(g382), .CK(CK) );
DFF_X2 U_g383 ( .D(g382), .Q(g383), .CK(CK) );
DFF_X2 U_g387 ( .D(g11506), .Q(g387), .CK(CK) );
DFF_X2 U_g394 ( .D(g387), .Q(g394), .CK(CK) );
DFF_X2 U_g395 ( .D(g11507), .Q(g395), .CK(CK) );
DFF_X2 U_g396 ( .D(g395), .Q(g396), .CK(CK) );
DFF_X2 U_g397 ( .D(g11508), .Q(g397), .CK(CK) );
DFF_X2 U_g324 ( .D(g397), .Q(g324), .CK(CK) );
DFF_X2 U_g325 ( .D(g13408), .Q(g325), .CK(CK) );
DFF_X2 U_g331 ( .D(g325), .Q(g331), .CK(CK) );
DFF_X2 U_g337 ( .D(g331), .Q(g337), .CK(CK) );
DFF_X2 U_g545 ( .D(g13419), .Q(g545), .CK(CK) );
DFF_X2 U_g551 ( .D(g545), .Q(g551), .CK(CK) );
DFF_X2 U_g550 ( .D(g551), .Q(g550), .CK(CK) );
DFF_X2 U_g554 ( .D(g23160), .Q(g554), .CK(CK) );
DFF_X2 U_g557 ( .D(g20556), .Q(g557), .CK(CK) );
DFF_X2 U_g510 ( .D(g20557), .Q(g510), .CK(CK) );
DFF_X2 U_g513 ( .D(g16467), .Q(g513), .CK(CK) );
DFF_X2 U_g523 ( .D(g513), .Q(g523), .CK(CK) );
DFF_X2 U_g524 ( .D(g523), .Q(g524), .CK(CK) );
DFF_X2 U_g564 ( .D(g11512), .Q(g564), .CK(CK) );
DFF_X2 U_g569 ( .D(g564), .Q(g569), .CK(CK) );
DFF_X2 U_g570 ( .D(g11515), .Q(g570), .CK(CK) );
DFF_X2 U_g571 ( .D(g570), .Q(g571), .CK(CK) );
DFF_X2 U_g572 ( .D(g11516), .Q(g572), .CK(CK) );
DFF_X2 U_g573 ( .D(g572), .Q(g573), .CK(CK) );
DFF_X2 U_g574 ( .D(g11517), .Q(g574), .CK(CK) );
DFF_X2 U_g565 ( .D(g574), .Q(g565), .CK(CK) );
DFF_X2 U_g566 ( .D(g11513), .Q(g566), .CK(CK) );
DFF_X2 U_g567 ( .D(g566), .Q(g567), .CK(CK) );
DFF_X2 U_g568 ( .D(g11514), .Q(g568), .CK(CK) );
DFF_X2 U_g489 ( .D(g568), .Q(g489), .CK(CK) );
DFF_X2 U_g474 ( .D(g13409), .Q(g474), .CK(CK) );
DFF_X2 U_g481 ( .D(g474), .Q(g481), .CK(CK) );
DFF_X2 U_g485 ( .D(g481), .Q(g485), .CK(CK) );
DFF_X2 U_g486 ( .D(g24292), .Q(g486), .CK(CK) );
DFF_X2 U_g487 ( .D(g24293), .Q(g487), .CK(CK) );
DFF_X2 U_g488 ( .D(g24294), .Q(g488), .CK(CK) );
DFF_X2 U_g455 ( .D(g25139), .Q(g455), .CK(CK) );
DFF_X2 U_g458 ( .D(g25131), .Q(g458), .CK(CK) );
DFF_X2 U_g461 ( .D(g25132), .Q(g461), .CK(CK) );
DFF_X2 U_g477 ( .D(g25136), .Q(g477), .CK(CK) );
DFF_X2 U_g478 ( .D(g25137), .Q(g478), .CK(CK) );
DFF_X2 U_g479 ( .D(g25138), .Q(g479), .CK(CK) );
DFF_X2 U_g480 ( .D(g24289), .Q(g480), .CK(CK) );
DFF_X2 U_g484 ( .D(g24290), .Q(g484), .CK(CK) );
DFF_X2 U_g464 ( .D(g24291), .Q(g464), .CK(CK) );
DFF_X2 U_g465 ( .D(g25133), .Q(g465), .CK(CK) );
DFF_X2 U_g468 ( .D(g25134), .Q(g468), .CK(CK) );
DFF_X2 U_g471 ( .D(g25135), .Q(g471), .CK(CK) );
DFF_X2 U_g528 ( .D(g16468), .Q(g528), .CK(CK) );
DFF_X2 U_g535 ( .D(g528), .Q(g535), .CK(CK) );
DFF_X2 U_g542 ( .D(g535), .Q(g542), .CK(CK) );
DFF_X2 U_g543 ( .D(g19021), .Q(g543), .CK(CK) );
DFF_X2 U_g544 ( .D(g543), .Q(g544), .CK(CK) );
DFF_X2 U_g548 ( .D(g23159), .Q(g548), .CK(CK) );
DFF_X2 U_g549 ( .D(g19022), .Q(g549), .CK(CK) );
DFF_X2 U_g499 ( .D(g549), .Q(g499), .CK(CK) );
DFF_X2 U_g558 ( .D(g19023), .Q(g558), .CK(CK) );
DFF_X2 U_g559 ( .D(g558), .Q(g559), .CK(CK) );
DFF_X2 U_g576 ( .D(g28219), .Q(g576), .CK(CK) );
DFF_X2 U_g577 ( .D(g28220), .Q(g577), .CK(CK) );
DFF_X2 U_g575 ( .D(g28221), .Q(g575), .CK(CK) );
DFF_X2 U_g579 ( .D(g28222), .Q(g579), .CK(CK) );
DFF_X2 U_g580 ( .D(g28223), .Q(g580), .CK(CK) );
DFF_X2 U_g578 ( .D(g28224), .Q(g578), .CK(CK) );
DFF_X2 U_g582 ( .D(g28225), .Q(g582), .CK(CK) );
DFF_X2 U_g583 ( .D(g28226), .Q(g583), .CK(CK) );
DFF_X2 U_g581 ( .D(g28227), .Q(g581), .CK(CK) );
DFF_X2 U_g585 ( .D(g28228), .Q(g585), .CK(CK) );
DFF_X2 U_g586 ( .D(g28229), .Q(g586), .CK(CK) );
DFF_X2 U_g584 ( .D(g28230), .Q(g584), .CK(CK) );
DFF_X2 U_g587 ( .D(g25985), .Q(g587), .CK(CK) );
DFF_X2 U_g590 ( .D(g25986), .Q(g590), .CK(CK) );
DFF_X2 U_g593 ( .D(g25987), .Q(g593), .CK(CK) );
DFF_X2 U_g596 ( .D(g25988), .Q(g596), .CK(CK) );
DFF_X2 U_g599 ( .D(g25989), .Q(g599), .CK(CK) );
DFF_X2 U_g602 ( .D(g25990), .Q(g602), .CK(CK) );
DFF_X2 U_g614 ( .D(g29135), .Q(g614), .CK(CK) );
DFF_X2 U_g617 ( .D(g29136), .Q(g617), .CK(CK) );
DFF_X2 U_g620 ( .D(g29137), .Q(g620), .CK(CK) );
DFF_X2 U_g605 ( .D(g29132), .Q(g605), .CK(CK) );
DFF_X2 U_g608 ( .D(g29133), .Q(g608), .CK(CK) );
DFF_X2 U_g611 ( .D(g29134), .Q(g611), .CK(CK) );
DFF_X2 U_g490 ( .D(g27194), .Q(g490), .CK(CK) );
DFF_X2 U_g493 ( .D(g27195), .Q(g493), .CK(CK) );
DFF_X2 U_g496 ( .D(g27196), .Q(g496), .CK(CK) );
DFF_X2 U_g506 ( .D(g8284), .Q(g506), .CK(CK) );
DFF_X2 U_g507 ( .D(g24295), .Q(g507), .CK(CK) );
DFF_X2 U_g508 ( .D(g19017), .Q(g508), .CK(CK) );
DFF_X2 U_g509 ( .D(g19018), .Q(g509), .CK(CK) );
DFF_X2 U_g514 ( .D(g19019), .Q(g514), .CK(CK) );
DFF_X2 U_g515 ( .D(g19020), .Q(g515), .CK(CK) );
DFF_X2 U_g516 ( .D(g23158), .Q(g516), .CK(CK) );
DFF_X2 U_g517 ( .D(g23157), .Q(g517), .CK(CK) );
DFF_X2 U_g518 ( .D(g23156), .Q(g518), .CK(CK) );
DFF_X2 U_g519 ( .D(g23155), .Q(g519), .CK(CK) );
DFF_X2 U_g520 ( .D(g23154), .Q(g520), .CK(CK) );
DFF_X2 U_g525 ( .D(g520), .Q(g525), .CK(CK) );
DFF_X2 U_g529 ( .D(g13410), .Q(g529), .CK(CK) );
DFF_X2 U_g530 ( .D(g13411), .Q(g530), .CK(CK) );
DFF_X2 U_g531 ( .D(g13412), .Q(g531), .CK(CK) );
DFF_X2 U_g532 ( .D(g13413), .Q(g532), .CK(CK) );
DFF_X2 U_g533 ( .D(g13414), .Q(g533), .CK(CK) );
DFF_X2 U_g534 ( .D(g13415), .Q(g534), .CK(CK) );
DFF_X2 U_g536 ( .D(g13416), .Q(g536), .CK(CK) );
DFF_X2 U_g537 ( .D(g13417), .Q(g537), .CK(CK) );
DFF_X2 U_g538 ( .D(g25984), .Q(g538), .CK(CK) );
DFF_X2 U_g541 ( .D(g13418), .Q(g541), .CK(CK) );
DFF_X2 U_g623 ( .D(g13420), .Q(g623), .CK(CK) );
DFF_X2 U_g626 ( .D(g623), .Q(g626), .CK(CK) );
DFF_X2 U_g629 ( .D(g626), .Q(g629), .CK(CK) );
DFF_X2 U_g630 ( .D(g20558), .Q(g630), .CK(CK) );
DFF_X2 U_g659 ( .D(g21943), .Q(g659), .CK(CK) );
DFF_X2 U_g640 ( .D(g23161), .Q(g640), .CK(CK) );
DFF_X2 U_g633 ( .D(g24296), .Q(g633), .CK(CK) );
DFF_X2 U_g653 ( .D(g25140), .Q(g653), .CK(CK) );
DFF_X2 U_g646 ( .D(g25991), .Q(g646), .CK(CK) );
DFF_X2 U_g660 ( .D(g26691), .Q(g660), .CK(CK) );
DFF_X2 U_g672 ( .D(g27197), .Q(g672), .CK(CK) );
DFF_X2 U_g666 ( .D(g27690), .Q(g666), .CK(CK) );
DFF_X2 U_g679 ( .D(g28231), .Q(g679), .CK(CK) );
DFF_X2 U_g686 ( .D(g28677), .Q(g686), .CK(CK) );
DFF_X2 U_g692 ( .D(g29138), .Q(g692), .CK(CK) );
DFF_X2 U_g699 ( .D(g23162), .Q(g699), .CK(CK) );
DFF_X2 U_g700 ( .D(g23163), .Q(g700), .CK(CK) );
DFF_X2 U_g698 ( .D(g23164), .Q(g698), .CK(CK) );
DFF_X2 U_g702 ( .D(g23165), .Q(g702), .CK(CK) );
DFF_X2 U_g703 ( .D(g23166), .Q(g703), .CK(CK) );
DFF_X2 U_g701 ( .D(g23167), .Q(g701), .CK(CK) );
DFF_X2 U_g705 ( .D(g23168), .Q(g705), .CK(CK) );
DFF_X2 U_g706 ( .D(g23169), .Q(g706), .CK(CK) );
DFF_X2 U_g704 ( .D(g23170), .Q(g704), .CK(CK) );
DFF_X2 U_g708 ( .D(g23171), .Q(g708), .CK(CK) );
DFF_X2 U_g709 ( .D(g23172), .Q(g709), .CK(CK) );
DFF_X2 U_g707 ( .D(g23173), .Q(g707), .CK(CK) );
DFF_X2 U_g711 ( .D(g23174), .Q(g711), .CK(CK) );
DFF_X2 U_g712 ( .D(g23175), .Q(g712), .CK(CK) );
DFF_X2 U_g710 ( .D(g23176), .Q(g710), .CK(CK) );
DFF_X2 U_g714 ( .D(g23177), .Q(g714), .CK(CK) );
DFF_X2 U_g715 ( .D(g23178), .Q(g715), .CK(CK) );
DFF_X2 U_g713 ( .D(g23179), .Q(g713), .CK(CK) );
DFF_X2 U_g717 ( .D(g23180), .Q(g717), .CK(CK) );
DFF_X2 U_g718 ( .D(g23181), .Q(g718), .CK(CK) );
DFF_X2 U_g716 ( .D(g23182), .Q(g716), .CK(CK) );
DFF_X2 U_g720 ( .D(g23183), .Q(g720), .CK(CK) );
DFF_X2 U_g721 ( .D(g23184), .Q(g721), .CK(CK) );
DFF_X2 U_g719 ( .D(g23185), .Q(g719), .CK(CK) );
DFF_X2 U_g723 ( .D(g23186), .Q(g723), .CK(CK) );
DFF_X2 U_g724 ( .D(g23187), .Q(g724), .CK(CK) );
DFF_X2 U_g722 ( .D(g23188), .Q(g722), .CK(CK) );
DFF_X2 U_g726 ( .D(g23189), .Q(g726), .CK(CK) );
DFF_X2 U_g727 ( .D(g23190), .Q(g727), .CK(CK) );
DFF_X2 U_g725 ( .D(g23191), .Q(g725), .CK(CK) );
DFF_X2 U_g729 ( .D(g23192), .Q(g729), .CK(CK) );
DFF_X2 U_g730 ( .D(g23193), .Q(g730), .CK(CK) );
DFF_X2 U_g728 ( .D(g23194), .Q(g728), .CK(CK) );
DFF_X2 U_g732 ( .D(g23195), .Q(g732), .CK(CK) );
DFF_X2 U_g733 ( .D(g23196), .Q(g733), .CK(CK) );
DFF_X2 U_g731 ( .D(g23197), .Q(g731), .CK(CK) );
DFF_X2 U_g735 ( .D(g26692), .Q(g735), .CK(CK) );
DFF_X2 U_g736 ( .D(g26693), .Q(g736), .CK(CK) );
DFF_X2 U_g734 ( .D(g26694), .Q(g734), .CK(CK) );
DFF_X2 U_g738 ( .D(g24297), .Q(g738), .CK(CK) );
DFF_X2 U_g739 ( .D(g24298), .Q(g739), .CK(CK) );
DFF_X2 U_g737 ( .D(g24299), .Q(g737), .CK(CK) );
DFF_X2 U_g826 ( .D(g13421), .Q(g826), .CK(CK) );
DFF_X2 U_g823 ( .D(g826), .Q(g823), .CK(CK) );
DFF_X2 U_g853 ( .D(g823), .Q(g853), .CK(CK) );
DFF_X2 U_g818 ( .D(g24300), .Q(g818), .CK(CK) );
DFF_X2 U_g819 ( .D(g24301), .Q(g819), .CK(CK) );
DFF_X2 U_g817 ( .D(g24302), .Q(g817), .CK(CK) );
DFF_X2 U_g821 ( .D(g24303), .Q(g821), .CK(CK) );
DFF_X2 U_g822 ( .D(g24304), .Q(g822), .CK(CK) );
DFF_X2 U_g820 ( .D(g24305), .Q(g820), .CK(CK) );
DFF_X2 U_g830 ( .D(g24306), .Q(g830), .CK(CK) );
DFF_X2 U_g831 ( .D(g24307), .Q(g831), .CK(CK) );
DFF_X2 U_g829 ( .D(g24308), .Q(g829), .CK(CK) );
DFF_X2 U_g833 ( .D(g24309), .Q(g833), .CK(CK) );
DFF_X2 U_g834 ( .D(g24310), .Q(g834), .CK(CK) );
DFF_X2 U_g832 ( .D(g24311), .Q(g832), .CK(CK) );
DFF_X2 U_g836 ( .D(g24312), .Q(g836), .CK(CK) );
DFF_X2 U_g837 ( .D(g24313), .Q(g837), .CK(CK) );
DFF_X2 U_g835 ( .D(g24314), .Q(g835), .CK(CK) );
DFF_X2 U_g839 ( .D(g24315), .Q(g839), .CK(CK) );
DFF_X2 U_g840 ( .D(g24316), .Q(g840), .CK(CK) );
DFF_X2 U_g838 ( .D(g24317), .Q(g838), .CK(CK) );
DFF_X2 U_g842 ( .D(g24318), .Q(g842), .CK(CK) );
DFF_X2 U_g843 ( .D(g24319), .Q(g843), .CK(CK) );
DFF_X2 U_g841 ( .D(g24320), .Q(g841), .CK(CK) );
DFF_X2 U_g845 ( .D(g24321), .Q(g845), .CK(CK) );
DFF_X2 U_g846 ( .D(g24322), .Q(g846), .CK(CK) );
DFF_X2 U_g844 ( .D(g24323), .Q(g844), .CK(CK) );
DFF_X2 U_g848 ( .D(g24324), .Q(g848), .CK(CK) );
DFF_X2 U_g849 ( .D(g24325), .Q(g849), .CK(CK) );
DFF_X2 U_g847 ( .D(g24326), .Q(g847), .CK(CK) );
DFF_X2 U_g851 ( .D(g24327), .Q(g851), .CK(CK) );
DFF_X2 U_g852 ( .D(g24328), .Q(g852), .CK(CK) );
DFF_X2 U_g850 ( .D(g24329), .Q(g850), .CK(CK) );
DFF_X2 U_g857 ( .D(g26696), .Q(g857), .CK(CK) );
DFF_X2 U_g858 ( .D(g26697), .Q(g858), .CK(CK) );
DFF_X2 U_g856 ( .D(g26698), .Q(g856), .CK(CK) );
DFF_X2 U_g860 ( .D(g26699), .Q(g860), .CK(CK) );
DFF_X2 U_g861 ( .D(g26700), .Q(g861), .CK(CK) );
DFF_X2 U_g859 ( .D(g26701), .Q(g859), .CK(CK) );
DFF_X2 U_g863 ( .D(g26702), .Q(g863), .CK(CK) );
DFF_X2 U_g864 ( .D(g26703), .Q(g864), .CK(CK) );
DFF_X2 U_g862 ( .D(g26704), .Q(g862), .CK(CK) );
DFF_X2 U_g866 ( .D(g26705), .Q(g866), .CK(CK) );
DFF_X2 U_g867 ( .D(g26706), .Q(g867), .CK(CK) );
DFF_X2 U_g865 ( .D(g26707), .Q(g865), .CK(CK) );
DFF_X2 U_g873 ( .D(g30521), .Q(g873), .CK(CK) );
DFF_X2 U_g876 ( .D(g30522), .Q(g876), .CK(CK) );
DFF_X2 U_g879 ( .D(g30523), .Q(g879), .CK(CK) );
DFF_X2 U_g918 ( .D(g30860), .Q(g918), .CK(CK) );
DFF_X2 U_g921 ( .D(g30861), .Q(g921), .CK(CK) );
DFF_X2 U_g924 ( .D(g30862), .Q(g924), .CK(CK) );
DFF_X2 U_g882 ( .D(g30854), .Q(g882), .CK(CK) );
DFF_X2 U_g885 ( .D(g30855), .Q(g885), .CK(CK) );
DFF_X2 U_g888 ( .D(g30856), .Q(g888), .CK(CK) );
DFF_X2 U_g927 ( .D(g30863), .Q(g927), .CK(CK) );
DFF_X2 U_g930 ( .D(g30864), .Q(g930), .CK(CK) );
DFF_X2 U_g933 ( .D(g30865), .Q(g933), .CK(CK) );
DFF_X2 U_g891 ( .D(g30524), .Q(g891), .CK(CK) );
DFF_X2 U_g894 ( .D(g30525), .Q(g894), .CK(CK) );
DFF_X2 U_g897 ( .D(g30526), .Q(g897), .CK(CK) );
DFF_X2 U_g936 ( .D(g30530), .Q(g936), .CK(CK) );
DFF_X2 U_g939 ( .D(g30531), .Q(g939), .CK(CK) );
DFF_X2 U_g942 ( .D(g30532), .Q(g942), .CK(CK) );
DFF_X2 U_g900 ( .D(g30527), .Q(g900), .CK(CK) );
DFF_X2 U_g903 ( .D(g30528), .Q(g903), .CK(CK) );
DFF_X2 U_g906 ( .D(g30529), .Q(g906), .CK(CK) );
DFF_X2 U_g945 ( .D(g30533), .Q(g945), .CK(CK) );
DFF_X2 U_g948 ( .D(g30534), .Q(g948), .CK(CK) );
DFF_X2 U_g951 ( .D(g30535), .Q(g951), .CK(CK) );
DFF_X2 U_g909 ( .D(g30857), .Q(g909), .CK(CK) );
DFF_X2 U_g912 ( .D(g30858), .Q(g912), .CK(CK) );
DFF_X2 U_g915 ( .D(g30859), .Q(g915), .CK(CK) );
DFF_X2 U_g954 ( .D(g30866), .Q(g954), .CK(CK) );
DFF_X2 U_g957 ( .D(g30867), .Q(g957), .CK(CK) );
DFF_X2 U_g960 ( .D(g30868), .Q(g960), .CK(CK) );
DFF_X2 U_g780 ( .D(g25992), .Q(g780), .CK(CK) );
DFF_X2 U_g776 ( .D(g26695), .Q(g776), .CK(CK) );
DFF_X2 U_g771 ( .D(g27198), .Q(g771), .CK(CK) );
DFF_X2 U_g767 ( .D(g27691), .Q(g767), .CK(CK) );
DFF_X2 U_g762 ( .D(g28232), .Q(g762), .CK(CK) );
DFF_X2 U_g758 ( .D(g28678), .Q(g758), .CK(CK) );
DFF_X2 U_g753 ( .D(g29139), .Q(g753), .CK(CK) );
DFF_X2 U_g749 ( .D(g29420), .Q(g749), .CK(CK) );
DFF_X2 U_g744 ( .D(g29634), .Q(g744), .CK(CK) );
DFF_X2 U_g740 ( .D(g29798), .Q(g740), .CK(CK) );
DFF_X2 U_g868 ( .D(g20559), .Q(g868), .CK(CK) );
DFF_X2 U_g870 ( .D(g868), .Q(g870), .CK(CK) );
DFF_X2 U_g869 ( .D(g870), .Q(g869), .CK(CK) );
DFF_X2 U_g963 ( .D(g13422), .Q(g963), .CK(CK) );
DFF_X2 U_g1092 ( .D(g963), .Q(g1092), .CK(CK) );
DFF_X2 U_g1088 ( .D(g1092), .Q(g1088), .CK(CK) );
DFF_X2 U_g996 ( .D(g11523), .Q(g996), .CK(CK) );
DFF_X2 U_g1041 ( .D(g28233), .Q(g1041), .CK(CK) );
DFF_X2 U_g1030 ( .D(g28234), .Q(g1030), .CK(CK) );
DFF_X2 U_g1033 ( .D(g28235), .Q(g1033), .CK(CK) );
DFF_X2 U_g1056 ( .D(g28236), .Q(g1056), .CK(CK) );
DFF_X2 U_g1045 ( .D(g28237), .Q(g1045), .CK(CK) );
DFF_X2 U_g1048 ( .D(g28238), .Q(g1048), .CK(CK) );
DFF_X2 U_g1071 ( .D(g28239), .Q(g1071), .CK(CK) );
DFF_X2 U_g1060 ( .D(g28240), .Q(g1060), .CK(CK) );
DFF_X2 U_g1063 ( .D(g28241), .Q(g1063), .CK(CK) );
DFF_X2 U_g1085 ( .D(g28242), .Q(g1085), .CK(CK) );
DFF_X2 U_g1075 ( .D(g28243), .Q(g1075), .CK(CK) );
DFF_X2 U_g1078 ( .D(g28244), .Q(g1078), .CK(CK) );
DFF_X2 U_g1095 ( .D(g29421), .Q(g1095), .CK(CK) );
DFF_X2 U_g1098 ( .D(g29422), .Q(g1098), .CK(CK) );
DFF_X2 U_g1101 ( .D(g29423), .Q(g1101), .CK(CK) );
DFF_X2 U_g1104 ( .D(g29638), .Q(g1104), .CK(CK) );
DFF_X2 U_g1107 ( .D(g29639), .Q(g1107), .CK(CK) );
DFF_X2 U_g1110 ( .D(g29640), .Q(g1110), .CK(CK) );
DFF_X2 U_g1114 ( .D(g29424), .Q(g1114), .CK(CK) );
DFF_X2 U_g1115 ( .D(g29425), .Q(g1115), .CK(CK) );
DFF_X2 U_g1113 ( .D(g29426), .Q(g1113), .CK(CK) );
DFF_X2 U_g1116 ( .D(g27692), .Q(g1116), .CK(CK) );
DFF_X2 U_g1119 ( .D(g27693), .Q(g1119), .CK(CK) );
DFF_X2 U_g1122 ( .D(g27694), .Q(g1122), .CK(CK) );
DFF_X2 U_g1125 ( .D(g27695), .Q(g1125), .CK(CK) );
DFF_X2 U_g1128 ( .D(g27696), .Q(g1128), .CK(CK) );
DFF_X2 U_g1131 ( .D(g27697), .Q(g1131), .CK(CK) );
DFF_X2 U_g1135 ( .D(g28679), .Q(g1135), .CK(CK) );
DFF_X2 U_g1136 ( .D(g28680), .Q(g1136), .CK(CK) );
DFF_X2 U_g1134 ( .D(g28681), .Q(g1134), .CK(CK) );
DFF_X2 U_g999 ( .D(g29799), .Q(g999), .CK(CK) );
DFF_X2 U_g1000 ( .D(g29800), .Q(g1000), .CK(CK) );
DFF_X2 U_g1001 ( .D(g29801), .Q(g1001), .CK(CK) );
DFF_X2 U_g1002 ( .D(g30869), .Q(g1002), .CK(CK) );
DFF_X2 U_g1003 ( .D(g30870), .Q(g1003), .CK(CK) );
DFF_X2 U_g1004 ( .D(g30871), .Q(g1004), .CK(CK) );
DFF_X2 U_g1005 ( .D(g30713), .Q(g1005), .CK(CK) );
DFF_X2 U_g1006 ( .D(g30714), .Q(g1006), .CK(CK) );
DFF_X2 U_g1007 ( .D(g30715), .Q(g1007), .CK(CK) );
DFF_X2 U_g1009 ( .D(g29635), .Q(g1009), .CK(CK) );
DFF_X2 U_g1010 ( .D(g29636), .Q(g1010), .CK(CK) );
DFF_X2 U_g1008 ( .D(g29637), .Q(g1008), .CK(CK) );
DFF_X2 U_g1090 ( .D(g27206), .Q(g1090), .CK(CK) );
DFF_X2 U_g1091 ( .D(g27207), .Q(g1091), .CK(CK) );
DFF_X2 U_g1089 ( .D(g27208), .Q(g1089), .CK(CK) );
DFF_X2 U_g1137 ( .D(g11536), .Q(g1137), .CK(CK) );
DFF_X2 U_g1138 ( .D(g1137), .Q(g1138), .CK(CK) );
DFF_X2 U_g1139 ( .D(g11537), .Q(g1139), .CK(CK) );
DFF_X2 U_g1140 ( .D(g1139), .Q(g1140), .CK(CK) );
DFF_X2 U_g1141 ( .D(g11538), .Q(g1141), .CK(CK) );
DFF_X2 U_g966 ( .D(g1141), .Q(g966), .CK(CK) );
DFF_X2 U_g967 ( .D(g11518), .Q(g967), .CK(CK) );
DFF_X2 U_g968 ( .D(g967), .Q(g968), .CK(CK) );
DFF_X2 U_g969 ( .D(g11519), .Q(g969), .CK(CK) );
DFF_X2 U_g970 ( .D(g969), .Q(g970), .CK(CK) );
DFF_X2 U_g971 ( .D(g11520), .Q(g971), .CK(CK) );
DFF_X2 U_g972 ( .D(g971), .Q(g972), .CK(CK) );
DFF_X2 U_g973 ( .D(g11521), .Q(g973), .CK(CK) );
DFF_X2 U_g974 ( .D(g973), .Q(g974), .CK(CK) );
DFF_X2 U_g975 ( .D(g11522), .Q(g975), .CK(CK) );
DFF_X2 U_g976 ( .D(g975), .Q(g976), .CK(CK) );
DFF_X2 U_g977 ( .D(g13423), .Q(g977), .CK(CK) );
DFF_X2 U_g978 ( .D(g977), .Q(g978), .CK(CK) );
DFF_X2 U_g986 ( .D(g19024), .Q(g986), .CK(CK) );
DFF_X2 U_g992 ( .D(g27200), .Q(g992), .CK(CK) );
DFF_X2 U_g995 ( .D(g27201), .Q(g995), .CK(CK) );
DFF_X2 U_g984 ( .D(g27202), .Q(g984), .CK(CK) );
DFF_X2 U_g983 ( .D(g27203), .Q(g983), .CK(CK) );
DFF_X2 U_g982 ( .D(g27204), .Q(g982), .CK(CK) );
DFF_X2 U_g981 ( .D(g27205), .Q(g981), .CK(CK) );
DFF_X2 U_g991 ( .D(g19028), .Q(g991), .CK(CK) );
DFF_X2 U_g990 ( .D(g19027), .Q(g990), .CK(CK) );
DFF_X2 U_g989 ( .D(g19026), .Q(g989), .CK(CK) );
DFF_X2 U_g988 ( .D(g19025), .Q(g988), .CK(CK) );
DFF_X2 U_g987 ( .D(g25141), .Q(g987), .CK(CK) );
DFF_X2 U_g985 ( .D(g27199), .Q(g985), .CK(CK) );
DFF_X2 U_g1029 ( .D(g11524), .Q(g1029), .CK(CK) );
DFF_X2 U_g1036 ( .D(g1029), .Q(g1036), .CK(CK) );
DFF_X2 U_g1037 ( .D(g11525), .Q(g1037), .CK(CK) );
DFF_X2 U_g1038 ( .D(g1037), .Q(g1038), .CK(CK) );
DFF_X2 U_g1039 ( .D(g11526), .Q(g1039), .CK(CK) );
DFF_X2 U_g1040 ( .D(g1039), .Q(g1040), .CK(CK) );
DFF_X2 U_g1044 ( .D(g11527), .Q(g1044), .CK(CK) );
DFF_X2 U_g1051 ( .D(g1044), .Q(g1051), .CK(CK) );
DFF_X2 U_g1052 ( .D(g11528), .Q(g1052), .CK(CK) );
DFF_X2 U_g1053 ( .D(g1052), .Q(g1053), .CK(CK) );
DFF_X2 U_g1054 ( .D(g11529), .Q(g1054), .CK(CK) );
DFF_X2 U_g1055 ( .D(g1054), .Q(g1055), .CK(CK) );
DFF_X2 U_g1059 ( .D(g11530), .Q(g1059), .CK(CK) );
DFF_X2 U_g1066 ( .D(g1059), .Q(g1066), .CK(CK) );
DFF_X2 U_g1067 ( .D(g11531), .Q(g1067), .CK(CK) );
DFF_X2 U_g1068 ( .D(g1067), .Q(g1068), .CK(CK) );
DFF_X2 U_g1069 ( .D(g11532), .Q(g1069), .CK(CK) );
DFF_X2 U_g1070 ( .D(g1069), .Q(g1070), .CK(CK) );
DFF_X2 U_g1074 ( .D(g11533), .Q(g1074), .CK(CK) );
DFF_X2 U_g1081 ( .D(g1074), .Q(g1081), .CK(CK) );
DFF_X2 U_g1082 ( .D(g11534), .Q(g1082), .CK(CK) );
DFF_X2 U_g1083 ( .D(g1082), .Q(g1083), .CK(CK) );
DFF_X2 U_g1084 ( .D(g11535), .Q(g1084), .CK(CK) );
DFF_X2 U_g1011 ( .D(g1084), .Q(g1011), .CK(CK) );
DFF_X2 U_g1012 ( .D(g13424), .Q(g1012), .CK(CK) );
DFF_X2 U_g1018 ( .D(g1012), .Q(g1018), .CK(CK) );
DFF_X2 U_g1024 ( .D(g1018), .Q(g1024), .CK(CK) );
DFF_X2 U_g1231 ( .D(g13435), .Q(g1231), .CK(CK) );
DFF_X2 U_g1237 ( .D(g1231), .Q(g1237), .CK(CK) );
DFF_X2 U_g1236 ( .D(g1237), .Q(g1236), .CK(CK) );
DFF_X2 U_g1240 ( .D(g23198), .Q(g1240), .CK(CK) );
DFF_X2 U_g1243 ( .D(g20560), .Q(g1243), .CK(CK) );
DFF_X2 U_g1196 ( .D(g20561), .Q(g1196), .CK(CK) );
DFF_X2 U_g1199 ( .D(g16469), .Q(g1199), .CK(CK) );
DFF_X2 U_g1209 ( .D(g1199), .Q(g1209), .CK(CK) );
DFF_X2 U_g1210 ( .D(g1209), .Q(g1210), .CK(CK) );
DFF_X2 U_g1250 ( .D(g11539), .Q(g1250), .CK(CK) );
DFF_X2 U_g1255 ( .D(g1250), .Q(g1255), .CK(CK) );
DFF_X2 U_g1256 ( .D(g11542), .Q(g1256), .CK(CK) );
DFF_X2 U_g1257 ( .D(g1256), .Q(g1257), .CK(CK) );
DFF_X2 U_g1258 ( .D(g11543), .Q(g1258), .CK(CK) );
DFF_X2 U_g1259 ( .D(g1258), .Q(g1259), .CK(CK) );
DFF_X2 U_g1260 ( .D(g11544), .Q(g1260), .CK(CK) );
DFF_X2 U_g1251 ( .D(g1260), .Q(g1251), .CK(CK) );
DFF_X2 U_g1252 ( .D(g11540), .Q(g1252), .CK(CK) );
DFF_X2 U_g1253 ( .D(g1252), .Q(g1253), .CK(CK) );
DFF_X2 U_g1254 ( .D(g11541), .Q(g1254), .CK(CK) );
DFF_X2 U_g1176 ( .D(g1254), .Q(g1176), .CK(CK) );
DFF_X2 U_g1161 ( .D(g13425), .Q(g1161), .CK(CK) );
DFF_X2 U_g1168 ( .D(g1161), .Q(g1168), .CK(CK) );
DFF_X2 U_g1172 ( .D(g1168), .Q(g1172), .CK(CK) );
DFF_X2 U_g1173 ( .D(g24333), .Q(g1173), .CK(CK) );
DFF_X2 U_g1174 ( .D(g24334), .Q(g1174), .CK(CK) );
DFF_X2 U_g1175 ( .D(g24335), .Q(g1175), .CK(CK) );
DFF_X2 U_g1142 ( .D(g25150), .Q(g1142), .CK(CK) );
DFF_X2 U_g1145 ( .D(g25142), .Q(g1145), .CK(CK) );
DFF_X2 U_g1148 ( .D(g25143), .Q(g1148), .CK(CK) );
DFF_X2 U_g1164 ( .D(g25147), .Q(g1164), .CK(CK) );
DFF_X2 U_g1165 ( .D(g25148), .Q(g1165), .CK(CK) );
DFF_X2 U_g1166 ( .D(g25149), .Q(g1166), .CK(CK) );
DFF_X2 U_g1167 ( .D(g24330), .Q(g1167), .CK(CK) );
DFF_X2 U_g1171 ( .D(g24331), .Q(g1171), .CK(CK) );
DFF_X2 U_g1151 ( .D(g24332), .Q(g1151), .CK(CK) );
DFF_X2 U_g1152 ( .D(g25144), .Q(g1152), .CK(CK) );
DFF_X2 U_g1155 ( .D(g25145), .Q(g1155), .CK(CK) );
DFF_X2 U_g1158 ( .D(g25146), .Q(g1158), .CK(CK) );
DFF_X2 U_g1214 ( .D(g16470), .Q(g1214), .CK(CK) );
DFF_X2 U_g1221 ( .D(g1214), .Q(g1221), .CK(CK) );
DFF_X2 U_g1228 ( .D(g1221), .Q(g1228), .CK(CK) );
DFF_X2 U_g1229 ( .D(g19033), .Q(g1229), .CK(CK) );
DFF_X2 U_g1230 ( .D(g1229), .Q(g1230), .CK(CK) );
DFF_X2 U_g1234 ( .D(g27217), .Q(g1234), .CK(CK) );
DFF_X2 U_g1235 ( .D(g19034), .Q(g1235), .CK(CK) );
DFF_X2 U_g1186 ( .D(g1235), .Q(g1186), .CK(CK) );
DFF_X2 U_g1244 ( .D(g19035), .Q(g1244), .CK(CK) );
DFF_X2 U_g1245 ( .D(g1244), .Q(g1245), .CK(CK) );
DFF_X2 U_g1262 ( .D(g28245), .Q(g1262), .CK(CK) );
DFF_X2 U_g1263 ( .D(g28246), .Q(g1263), .CK(CK) );
DFF_X2 U_g1261 ( .D(g28247), .Q(g1261), .CK(CK) );
DFF_X2 U_g1265 ( .D(g28248), .Q(g1265), .CK(CK) );
DFF_X2 U_g1266 ( .D(g28249), .Q(g1266), .CK(CK) );
DFF_X2 U_g1264 ( .D(g28250), .Q(g1264), .CK(CK) );
DFF_X2 U_g1268 ( .D(g28251), .Q(g1268), .CK(CK) );
DFF_X2 U_g1269 ( .D(g28252), .Q(g1269), .CK(CK) );
DFF_X2 U_g1267 ( .D(g28253), .Q(g1267), .CK(CK) );
DFF_X2 U_g1271 ( .D(g28254), .Q(g1271), .CK(CK) );
DFF_X2 U_g1272 ( .D(g28255), .Q(g1272), .CK(CK) );
DFF_X2 U_g1270 ( .D(g28256), .Q(g1270), .CK(CK) );
DFF_X2 U_g1273 ( .D(g25994), .Q(g1273), .CK(CK) );
DFF_X2 U_g1276 ( .D(g25995), .Q(g1276), .CK(CK) );
DFF_X2 U_g1279 ( .D(g25996), .Q(g1279), .CK(CK) );
DFF_X2 U_g1282 ( .D(g25997), .Q(g1282), .CK(CK) );
DFF_X2 U_g1285 ( .D(g25998), .Q(g1285), .CK(CK) );
DFF_X2 U_g1288 ( .D(g25999), .Q(g1288), .CK(CK) );
DFF_X2 U_g1300 ( .D(g29143), .Q(g1300), .CK(CK) );
DFF_X2 U_g1303 ( .D(g29144), .Q(g1303), .CK(CK) );
DFF_X2 U_g1306 ( .D(g29145), .Q(g1306), .CK(CK) );
DFF_X2 U_g1291 ( .D(g29140), .Q(g1291), .CK(CK) );
DFF_X2 U_g1294 ( .D(g29141), .Q(g1294), .CK(CK) );
DFF_X2 U_g1297 ( .D(g29142), .Q(g1297), .CK(CK) );
DFF_X2 U_g1177 ( .D(g27209), .Q(g1177), .CK(CK) );
DFF_X2 U_g1180 ( .D(g27210), .Q(g1180), .CK(CK) );
DFF_X2 U_g1183 ( .D(g27211), .Q(g1183), .CK(CK) );
DFF_X2 U_g1192 ( .D(g8293), .Q(g1192), .CK(CK) );
DFF_X2 U_g1193 ( .D(g24336), .Q(g1193), .CK(CK) );
DFF_X2 U_g1194 ( .D(g19029), .Q(g1194), .CK(CK) );
DFF_X2 U_g1195 ( .D(g19030), .Q(g1195), .CK(CK) );
DFF_X2 U_g1200 ( .D(g19031), .Q(g1200), .CK(CK) );
DFF_X2 U_g1201 ( .D(g19032), .Q(g1201), .CK(CK) );
DFF_X2 U_g1202 ( .D(g27216), .Q(g1202), .CK(CK) );
DFF_X2 U_g1203 ( .D(g27215), .Q(g1203), .CK(CK) );
DFF_X2 U_g1204 ( .D(g27214), .Q(g1204), .CK(CK) );
DFF_X2 U_g1205 ( .D(g27213), .Q(g1205), .CK(CK) );
DFF_X2 U_g1206 ( .D(g27212), .Q(g1206), .CK(CK) );
DFF_X2 U_g1211 ( .D(g1206), .Q(g1211), .CK(CK) );
DFF_X2 U_g1215 ( .D(g13426), .Q(g1215), .CK(CK) );
DFF_X2 U_g1216 ( .D(g13427), .Q(g1216), .CK(CK) );
DFF_X2 U_g1217 ( .D(g13428), .Q(g1217), .CK(CK) );
DFF_X2 U_g1218 ( .D(g13429), .Q(g1218), .CK(CK) );
DFF_X2 U_g1219 ( .D(g13430), .Q(g1219), .CK(CK) );
DFF_X2 U_g1220 ( .D(g13431), .Q(g1220), .CK(CK) );
DFF_X2 U_g1222 ( .D(g13432), .Q(g1222), .CK(CK) );
DFF_X2 U_g1223 ( .D(g13433), .Q(g1223), .CK(CK) );
DFF_X2 U_g1224 ( .D(g25993), .Q(g1224), .CK(CK) );
DFF_X2 U_g1227 ( .D(g13434), .Q(g1227), .CK(CK) );
DFF_X2 U_g1309 ( .D(g13436), .Q(g1309), .CK(CK) );
DFF_X2 U_g1312 ( .D(g1309), .Q(g1312), .CK(CK) );
DFF_X2 U_g1315 ( .D(g1312), .Q(g1315), .CK(CK) );
DFF_X2 U_g1316 ( .D(g20562), .Q(g1316), .CK(CK) );
DFF_X2 U_g1345 ( .D(g21944), .Q(g1345), .CK(CK) );
DFF_X2 U_g1326 ( .D(g23199), .Q(g1326), .CK(CK) );
DFF_X2 U_g1319 ( .D(g24337), .Q(g1319), .CK(CK) );
DFF_X2 U_g1339 ( .D(g25151), .Q(g1339), .CK(CK) );
DFF_X2 U_g1332 ( .D(g26000), .Q(g1332), .CK(CK) );
DFF_X2 U_g1346 ( .D(g26708), .Q(g1346), .CK(CK) );
DFF_X2 U_g1358 ( .D(g27218), .Q(g1358), .CK(CK) );
DFF_X2 U_g1352 ( .D(g27698), .Q(g1352), .CK(CK) );
DFF_X2 U_g1365 ( .D(g28257), .Q(g1365), .CK(CK) );
DFF_X2 U_g1372 ( .D(g28682), .Q(g1372), .CK(CK) );
DFF_X2 U_g1378 ( .D(g29146), .Q(g1378), .CK(CK) );
DFF_X2 U_g1385 ( .D(g23200), .Q(g1385), .CK(CK) );
DFF_X2 U_g1386 ( .D(g23201), .Q(g1386), .CK(CK) );
DFF_X2 U_g1384 ( .D(g23202), .Q(g1384), .CK(CK) );
DFF_X2 U_g1388 ( .D(g23203), .Q(g1388), .CK(CK) );
DFF_X2 U_g1389 ( .D(g23204), .Q(g1389), .CK(CK) );
DFF_X2 U_g1387 ( .D(g23205), .Q(g1387), .CK(CK) );
DFF_X2 U_g1391 ( .D(g23206), .Q(g1391), .CK(CK) );
DFF_X2 U_g1392 ( .D(g23207), .Q(g1392), .CK(CK) );
DFF_X2 U_g1390 ( .D(g23208), .Q(g1390), .CK(CK) );
DFF_X2 U_g1394 ( .D(g23209), .Q(g1394), .CK(CK) );
DFF_X2 U_g1395 ( .D(g23210), .Q(g1395), .CK(CK) );
DFF_X2 U_g1393 ( .D(g23211), .Q(g1393), .CK(CK) );
DFF_X2 U_g1397 ( .D(g23212), .Q(g1397), .CK(CK) );
DFF_X2 U_g1398 ( .D(g23213), .Q(g1398), .CK(CK) );
DFF_X2 U_g1396 ( .D(g23214), .Q(g1396), .CK(CK) );
DFF_X2 U_g1400 ( .D(g23215), .Q(g1400), .CK(CK) );
DFF_X2 U_g1401 ( .D(g23216), .Q(g1401), .CK(CK) );
DFF_X2 U_g1399 ( .D(g23217), .Q(g1399), .CK(CK) );
DFF_X2 U_g1403 ( .D(g23218), .Q(g1403), .CK(CK) );
DFF_X2 U_g1404 ( .D(g23219), .Q(g1404), .CK(CK) );
DFF_X2 U_g1402 ( .D(g23220), .Q(g1402), .CK(CK) );
DFF_X2 U_g1406 ( .D(g23221), .Q(g1406), .CK(CK) );
DFF_X2 U_g1407 ( .D(g23222), .Q(g1407), .CK(CK) );
DFF_X2 U_g1405 ( .D(g23223), .Q(g1405), .CK(CK) );
DFF_X2 U_g1409 ( .D(g23224), .Q(g1409), .CK(CK) );
DFF_X2 U_g1410 ( .D(g23225), .Q(g1410), .CK(CK) );
DFF_X2 U_g1408 ( .D(g23226), .Q(g1408), .CK(CK) );
DFF_X2 U_g1412 ( .D(g23227), .Q(g1412), .CK(CK) );
DFF_X2 U_g1413 ( .D(g23228), .Q(g1413), .CK(CK) );
DFF_X2 U_g1411 ( .D(g23229), .Q(g1411), .CK(CK) );
DFF_X2 U_g1415 ( .D(g23230), .Q(g1415), .CK(CK) );
DFF_X2 U_g1416 ( .D(g23231), .Q(g1416), .CK(CK) );
DFF_X2 U_g1414 ( .D(g23232), .Q(g1414), .CK(CK) );
DFF_X2 U_g1418 ( .D(g23233), .Q(g1418), .CK(CK) );
DFF_X2 U_g1419 ( .D(g23234), .Q(g1419), .CK(CK) );
DFF_X2 U_g1417 ( .D(g23235), .Q(g1417), .CK(CK) );
DFF_X2 U_g1421 ( .D(g26709), .Q(g1421), .CK(CK) );
DFF_X2 U_g1422 ( .D(g26710), .Q(g1422), .CK(CK) );
DFF_X2 U_g1420 ( .D(g26711), .Q(g1420), .CK(CK) );
DFF_X2 U_g1424 ( .D(g24338), .Q(g1424), .CK(CK) );
DFF_X2 U_g1425 ( .D(g24339), .Q(g1425), .CK(CK) );
DFF_X2 U_g1423 ( .D(g24340), .Q(g1423), .CK(CK) );
DFF_X2 U_g1520 ( .D(g13437), .Q(g1520), .CK(CK) );
DFF_X2 U_g1517 ( .D(g1520), .Q(g1517), .CK(CK) );
DFF_X2 U_g1547 ( .D(g1517), .Q(g1547), .CK(CK) );
DFF_X2 U_g1512 ( .D(g24341), .Q(g1512), .CK(CK) );
DFF_X2 U_g1513 ( .D(g24342), .Q(g1513), .CK(CK) );
DFF_X2 U_g1511 ( .D(g24343), .Q(g1511), .CK(CK) );
DFF_X2 U_g1515 ( .D(g24344), .Q(g1515), .CK(CK) );
DFF_X2 U_g1516 ( .D(g24345), .Q(g1516), .CK(CK) );
DFF_X2 U_g1514 ( .D(g24346), .Q(g1514), .CK(CK) );
DFF_X2 U_g1524 ( .D(g24347), .Q(g1524), .CK(CK) );
DFF_X2 U_g1525 ( .D(g24348), .Q(g1525), .CK(CK) );
DFF_X2 U_g1523 ( .D(g24349), .Q(g1523), .CK(CK) );
DFF_X2 U_g1527 ( .D(g24350), .Q(g1527), .CK(CK) );
DFF_X2 U_g1528 ( .D(g24351), .Q(g1528), .CK(CK) );
DFF_X2 U_g1526 ( .D(g24352), .Q(g1526), .CK(CK) );
DFF_X2 U_g1530 ( .D(g24353), .Q(g1530), .CK(CK) );
DFF_X2 U_g1531 ( .D(g24354), .Q(g1531), .CK(CK) );
DFF_X2 U_g1529 ( .D(g24355), .Q(g1529), .CK(CK) );
DFF_X2 U_g1533 ( .D(g24356), .Q(g1533), .CK(CK) );
DFF_X2 U_g1534 ( .D(g24357), .Q(g1534), .CK(CK) );
DFF_X2 U_g1532 ( .D(g24358), .Q(g1532), .CK(CK) );
DFF_X2 U_g1536 ( .D(g24359), .Q(g1536), .CK(CK) );
DFF_X2 U_g1537 ( .D(g24360), .Q(g1537), .CK(CK) );
DFF_X2 U_g1535 ( .D(g24361), .Q(g1535), .CK(CK) );
DFF_X2 U_g1539 ( .D(g24362), .Q(g1539), .CK(CK) );
DFF_X2 U_g1540 ( .D(g24363), .Q(g1540), .CK(CK) );
DFF_X2 U_g1538 ( .D(g24364), .Q(g1538), .CK(CK) );
DFF_X2 U_g1542 ( .D(g24365), .Q(g1542), .CK(CK) );
DFF_X2 U_g1543 ( .D(g24366), .Q(g1543), .CK(CK) );
DFF_X2 U_g1541 ( .D(g24367), .Q(g1541), .CK(CK) );
DFF_X2 U_g1545 ( .D(g24368), .Q(g1545), .CK(CK) );
DFF_X2 U_g1546 ( .D(g24369), .Q(g1546), .CK(CK) );
DFF_X2 U_g1544 ( .D(g24370), .Q(g1544), .CK(CK) );
DFF_X2 U_g1551 ( .D(g26713), .Q(g1551), .CK(CK) );
DFF_X2 U_g1552 ( .D(g26714), .Q(g1552), .CK(CK) );
DFF_X2 U_g1550 ( .D(g26715), .Q(g1550), .CK(CK) );
DFF_X2 U_g1554 ( .D(g26716), .Q(g1554), .CK(CK) );
DFF_X2 U_g1555 ( .D(g26717), .Q(g1555), .CK(CK) );
DFF_X2 U_g1553 ( .D(g26718), .Q(g1553), .CK(CK) );
DFF_X2 U_g1557 ( .D(g26719), .Q(g1557), .CK(CK) );
DFF_X2 U_g1558 ( .D(g26720), .Q(g1558), .CK(CK) );
DFF_X2 U_g1556 ( .D(g26721), .Q(g1556), .CK(CK) );
DFF_X2 U_g1560 ( .D(g26722), .Q(g1560), .CK(CK) );
DFF_X2 U_g1561 ( .D(g26723), .Q(g1561), .CK(CK) );
DFF_X2 U_g1559 ( .D(g26724), .Q(g1559), .CK(CK) );
DFF_X2 U_g1567 ( .D(g30536), .Q(g1567), .CK(CK) );
DFF_X2 U_g1570 ( .D(g30537), .Q(g1570), .CK(CK) );
DFF_X2 U_g1573 ( .D(g30538), .Q(g1573), .CK(CK) );
DFF_X2 U_g1612 ( .D(g30878), .Q(g1612), .CK(CK) );
DFF_X2 U_g1615 ( .D(g30879), .Q(g1615), .CK(CK) );
DFF_X2 U_g1618 ( .D(g30880), .Q(g1618), .CK(CK) );
DFF_X2 U_g1576 ( .D(g30872), .Q(g1576), .CK(CK) );
DFF_X2 U_g1579 ( .D(g30873), .Q(g1579), .CK(CK) );
DFF_X2 U_g1582 ( .D(g30874), .Q(g1582), .CK(CK) );
DFF_X2 U_g1621 ( .D(g30881), .Q(g1621), .CK(CK) );
DFF_X2 U_g1624 ( .D(g30882), .Q(g1624), .CK(CK) );
DFF_X2 U_g1627 ( .D(g30883), .Q(g1627), .CK(CK) );
DFF_X2 U_g1585 ( .D(g30539), .Q(g1585), .CK(CK) );
DFF_X2 U_g1588 ( .D(g30540), .Q(g1588), .CK(CK) );
DFF_X2 U_g1591 ( .D(g30541), .Q(g1591), .CK(CK) );
DFF_X2 U_g1630 ( .D(g30545), .Q(g1630), .CK(CK) );
DFF_X2 U_g1633 ( .D(g30546), .Q(g1633), .CK(CK) );
DFF_X2 U_g1636 ( .D(g30547), .Q(g1636), .CK(CK) );
DFF_X2 U_g1594 ( .D(g30542), .Q(g1594), .CK(CK) );
DFF_X2 U_g1597 ( .D(g30543), .Q(g1597), .CK(CK) );
DFF_X2 U_g1600 ( .D(g30544), .Q(g1600), .CK(CK) );
DFF_X2 U_g1639 ( .D(g30548), .Q(g1639), .CK(CK) );
DFF_X2 U_g1642 ( .D(g30549), .Q(g1642), .CK(CK) );
DFF_X2 U_g1645 ( .D(g30550), .Q(g1645), .CK(CK) );
DFF_X2 U_g1603 ( .D(g30875), .Q(g1603), .CK(CK) );
DFF_X2 U_g1606 ( .D(g30876), .Q(g1606), .CK(CK) );
DFF_X2 U_g1609 ( .D(g30877), .Q(g1609), .CK(CK) );
DFF_X2 U_g1648 ( .D(g30884), .Q(g1648), .CK(CK) );
DFF_X2 U_g1651 ( .D(g30885), .Q(g1651), .CK(CK) );
DFF_X2 U_g1654 ( .D(g30886), .Q(g1654), .CK(CK) );
DFF_X2 U_g1466 ( .D(g26001), .Q(g1466), .CK(CK) );
DFF_X2 U_g1462 ( .D(g26712), .Q(g1462), .CK(CK) );
DFF_X2 U_g1457 ( .D(g27219), .Q(g1457), .CK(CK) );
DFF_X2 U_g1453 ( .D(g27699), .Q(g1453), .CK(CK) );
DFF_X2 U_g1448 ( .D(g28258), .Q(g1448), .CK(CK) );
DFF_X2 U_g1444 ( .D(g28683), .Q(g1444), .CK(CK) );
DFF_X2 U_g1439 ( .D(g29147), .Q(g1439), .CK(CK) );
DFF_X2 U_g1435 ( .D(g29427), .Q(g1435), .CK(CK) );
DFF_X2 U_g1430 ( .D(g29641), .Q(g1430), .CK(CK) );
DFF_X2 U_g1426 ( .D(g29802), .Q(g1426), .CK(CK) );
DFF_X2 U_g1562 ( .D(g20563), .Q(g1562), .CK(CK) );
DFF_X2 U_g1564 ( .D(g1562), .Q(g1564), .CK(CK) );
DFF_X2 U_g1563 ( .D(g1564), .Q(g1563), .CK(CK) );
DFF_X2 U_g1657 ( .D(g13438), .Q(g1657), .CK(CK) );
DFF_X2 U_g1786 ( .D(g1657), .Q(g1786), .CK(CK) );
DFF_X2 U_g1782 ( .D(g1786), .Q(g1782), .CK(CK) );
DFF_X2 U_g1690 ( .D(g11550), .Q(g1690), .CK(CK) );
DFF_X2 U_g1735 ( .D(g28259), .Q(g1735), .CK(CK) );
DFF_X2 U_g1724 ( .D(g28260), .Q(g1724), .CK(CK) );
DFF_X2 U_g1727 ( .D(g28261), .Q(g1727), .CK(CK) );
DFF_X2 U_g1750 ( .D(g28262), .Q(g1750), .CK(CK) );
DFF_X2 U_g1739 ( .D(g28263), .Q(g1739), .CK(CK) );
DFF_X2 U_g1742 ( .D(g28264), .Q(g1742), .CK(CK) );
DFF_X2 U_g1765 ( .D(g28265), .Q(g1765), .CK(CK) );
DFF_X2 U_g1754 ( .D(g28266), .Q(g1754), .CK(CK) );
DFF_X2 U_g1757 ( .D(g28267), .Q(g1757), .CK(CK) );
DFF_X2 U_g1779 ( .D(g28268), .Q(g1779), .CK(CK) );
DFF_X2 U_g1769 ( .D(g28269), .Q(g1769), .CK(CK) );
DFF_X2 U_g1772 ( .D(g28270), .Q(g1772), .CK(CK) );
DFF_X2 U_g1789 ( .D(g29434), .Q(g1789), .CK(CK) );
DFF_X2 U_g1792 ( .D(g29435), .Q(g1792), .CK(CK) );
DFF_X2 U_g1795 ( .D(g29436), .Q(g1795), .CK(CK) );
DFF_X2 U_g1798 ( .D(g29645), .Q(g1798), .CK(CK) );
DFF_X2 U_g1801 ( .D(g29646), .Q(g1801), .CK(CK) );
DFF_X2 U_g1804 ( .D(g29647), .Q(g1804), .CK(CK) );
DFF_X2 U_g1808 ( .D(g29437), .Q(g1808), .CK(CK) );
DFF_X2 U_g1809 ( .D(g29438), .Q(g1809), .CK(CK) );
DFF_X2 U_g1807 ( .D(g29439), .Q(g1807), .CK(CK) );
DFF_X2 U_g1810 ( .D(g27700), .Q(g1810), .CK(CK) );
DFF_X2 U_g1813 ( .D(g27701), .Q(g1813), .CK(CK) );
DFF_X2 U_g1816 ( .D(g27702), .Q(g1816), .CK(CK) );
DFF_X2 U_g1819 ( .D(g27703), .Q(g1819), .CK(CK) );
DFF_X2 U_g1822 ( .D(g27704), .Q(g1822), .CK(CK) );
DFF_X2 U_g1825 ( .D(g27705), .Q(g1825), .CK(CK) );
DFF_X2 U_g1829 ( .D(g28684), .Q(g1829), .CK(CK) );
DFF_X2 U_g1830 ( .D(g28685), .Q(g1830), .CK(CK) );
DFF_X2 U_g1828 ( .D(g28686), .Q(g1828), .CK(CK) );
DFF_X2 U_g1693 ( .D(g29803), .Q(g1693), .CK(CK) );
DFF_X2 U_g1694 ( .D(g29804), .Q(g1694), .CK(CK) );
DFF_X2 U_g1695 ( .D(g29805), .Q(g1695), .CK(CK) );
DFF_X2 U_g1696 ( .D(g30887), .Q(g1696), .CK(CK) );
DFF_X2 U_g1697 ( .D(g30888), .Q(g1697), .CK(CK) );
DFF_X2 U_g1698 ( .D(g30889), .Q(g1698), .CK(CK) );
DFF_X2 U_g1699 ( .D(g30716), .Q(g1699), .CK(CK) );
DFF_X2 U_g1700 ( .D(g30717), .Q(g1700), .CK(CK) );
DFF_X2 U_g1701 ( .D(g30718), .Q(g1701), .CK(CK) );
DFF_X2 U_g1703 ( .D(g29642), .Q(g1703), .CK(CK) );
DFF_X2 U_g1704 ( .D(g29643), .Q(g1704), .CK(CK) );
DFF_X2 U_g1702 ( .D(g29644), .Q(g1702), .CK(CK) );
DFF_X2 U_g1784 ( .D(g27221), .Q(g1784), .CK(CK) );
DFF_X2 U_g1785 ( .D(g27222), .Q(g1785), .CK(CK) );
DFF_X2 U_g1783 ( .D(g27223), .Q(g1783), .CK(CK) );
DFF_X2 U_g1831 ( .D(g11563), .Q(g1831), .CK(CK) );
DFF_X2 U_g1832 ( .D(g1831), .Q(g1832), .CK(CK) );
DFF_X2 U_g1833 ( .D(g11564), .Q(g1833), .CK(CK) );
DFF_X2 U_g1834 ( .D(g1833), .Q(g1834), .CK(CK) );
DFF_X2 U_g1835 ( .D(g11565), .Q(g1835), .CK(CK) );
DFF_X2 U_g1660 ( .D(g1835), .Q(g1660), .CK(CK) );
DFF_X2 U_g1661 ( .D(g11545), .Q(g1661), .CK(CK) );
DFF_X2 U_g1662 ( .D(g1661), .Q(g1662), .CK(CK) );
DFF_X2 U_g1663 ( .D(g11546), .Q(g1663), .CK(CK) );
DFF_X2 U_g1664 ( .D(g1663), .Q(g1664), .CK(CK) );
DFF_X2 U_g1665 ( .D(g11547), .Q(g1665), .CK(CK) );
DFF_X2 U_g1666 ( .D(g1665), .Q(g1666), .CK(CK) );
DFF_X2 U_g1667 ( .D(g11548), .Q(g1667), .CK(CK) );
DFF_X2 U_g1668 ( .D(g1667), .Q(g1668), .CK(CK) );
DFF_X2 U_g1669 ( .D(g11549), .Q(g1669), .CK(CK) );
DFF_X2 U_g1670 ( .D(g1669), .Q(g1670), .CK(CK) );
DFF_X2 U_g1671 ( .D(g13439), .Q(g1671), .CK(CK) );
DFF_X2 U_g1672 ( .D(g1671), .Q(g1672), .CK(CK) );
DFF_X2 U_g1680 ( .D(g19036), .Q(g1680), .CK(CK) );
DFF_X2 U_g1686 ( .D(g29428), .Q(g1686), .CK(CK) );
DFF_X2 U_g1689 ( .D(g29429), .Q(g1689), .CK(CK) );
DFF_X2 U_g1678 ( .D(g29430), .Q(g1678), .CK(CK) );
DFF_X2 U_g1677 ( .D(g29431), .Q(g1677), .CK(CK) );
DFF_X2 U_g1676 ( .D(g29432), .Q(g1676), .CK(CK) );
DFF_X2 U_g1675 ( .D(g29433), .Q(g1675), .CK(CK) );
DFF_X2 U_g1685 ( .D(g19040), .Q(g1685), .CK(CK) );
DFF_X2 U_g1684 ( .D(g19039), .Q(g1684), .CK(CK) );
DFF_X2 U_g1683 ( .D(g19038), .Q(g1683), .CK(CK) );
DFF_X2 U_g1682 ( .D(g19037), .Q(g1682), .CK(CK) );
DFF_X2 U_g1681 ( .D(g25152), .Q(g1681), .CK(CK) );
DFF_X2 U_g1679 ( .D(g27220), .Q(g1679), .CK(CK) );
DFF_X2 U_g1723 ( .D(g11551), .Q(g1723), .CK(CK) );
DFF_X2 U_g1730 ( .D(g1723), .Q(g1730), .CK(CK) );
DFF_X2 U_g1731 ( .D(g11552), .Q(g1731), .CK(CK) );
DFF_X2 U_g1732 ( .D(g1731), .Q(g1732), .CK(CK) );
DFF_X2 U_g1733 ( .D(g11553), .Q(g1733), .CK(CK) );
DFF_X2 U_g1734 ( .D(g1733), .Q(g1734), .CK(CK) );
DFF_X2 U_g1738 ( .D(g11554), .Q(g1738), .CK(CK) );
DFF_X2 U_g1745 ( .D(g1738), .Q(g1745), .CK(CK) );
DFF_X2 U_g1746 ( .D(g11555), .Q(g1746), .CK(CK) );
DFF_X2 U_g1747 ( .D(g1746), .Q(g1747), .CK(CK) );
DFF_X2 U_g1748 ( .D(g11556), .Q(g1748), .CK(CK) );
DFF_X2 U_g1749 ( .D(g1748), .Q(g1749), .CK(CK) );
DFF_X2 U_g1753 ( .D(g11557), .Q(g1753), .CK(CK) );
DFF_X2 U_g1760 ( .D(g1753), .Q(g1760), .CK(CK) );
DFF_X2 U_g1761 ( .D(g11558), .Q(g1761), .CK(CK) );
DFF_X2 U_g1762 ( .D(g1761), .Q(g1762), .CK(CK) );
DFF_X2 U_g1763 ( .D(g11559), .Q(g1763), .CK(CK) );
DFF_X2 U_g1764 ( .D(g1763), .Q(g1764), .CK(CK) );
DFF_X2 U_g1768 ( .D(g11560), .Q(g1768), .CK(CK) );
DFF_X2 U_g1775 ( .D(g1768), .Q(g1775), .CK(CK) );
DFF_X2 U_g1776 ( .D(g11561), .Q(g1776), .CK(CK) );
DFF_X2 U_g1777 ( .D(g1776), .Q(g1777), .CK(CK) );
DFF_X2 U_g1778 ( .D(g11562), .Q(g1778), .CK(CK) );
DFF_X2 U_g1705 ( .D(g1778), .Q(g1705), .CK(CK) );
DFF_X2 U_g1706 ( .D(g13440), .Q(g1706), .CK(CK) );
DFF_X2 U_g1712 ( .D(g1706), .Q(g1712), .CK(CK) );
DFF_X2 U_g1718 ( .D(g1712), .Q(g1718), .CK(CK) );
DFF_X2 U_g1925 ( .D(g13451), .Q(g1925), .CK(CK) );
DFF_X2 U_g1931 ( .D(g1925), .Q(g1931), .CK(CK) );
DFF_X2 U_g1930 ( .D(g1931), .Q(g1930), .CK(CK) );
DFF_X2 U_g1934 ( .D(g23236), .Q(g1934), .CK(CK) );
DFF_X2 U_g1937 ( .D(g20564), .Q(g1937), .CK(CK) );
DFF_X2 U_g1890 ( .D(g20565), .Q(g1890), .CK(CK) );
DFF_X2 U_g1893 ( .D(g16471), .Q(g1893), .CK(CK) );
DFF_X2 U_g1903 ( .D(g1893), .Q(g1903), .CK(CK) );
DFF_X2 U_g1904 ( .D(g1903), .Q(g1904), .CK(CK) );
DFF_X2 U_g1944 ( .D(g11566), .Q(g1944), .CK(CK) );
DFF_X2 U_g1949 ( .D(g1944), .Q(g1949), .CK(CK) );
DFF_X2 U_g1950 ( .D(g11569), .Q(g1950), .CK(CK) );
DFF_X2 U_g1951 ( .D(g1950), .Q(g1951), .CK(CK) );
DFF_X2 U_g1952 ( .D(g11570), .Q(g1952), .CK(CK) );
DFF_X2 U_g1953 ( .D(g1952), .Q(g1953), .CK(CK) );
DFF_X2 U_g1954 ( .D(g11571), .Q(g1954), .CK(CK) );
DFF_X2 U_g1945 ( .D(g1954), .Q(g1945), .CK(CK) );
DFF_X2 U_g1946 ( .D(g11567), .Q(g1946), .CK(CK) );
DFF_X2 U_g1947 ( .D(g1946), .Q(g1947), .CK(CK) );
DFF_X2 U_g1948 ( .D(g11568), .Q(g1948), .CK(CK) );
DFF_X2 U_g1870 ( .D(g1948), .Q(g1870), .CK(CK) );
DFF_X2 U_g1855 ( .D(g13441), .Q(g1855), .CK(CK) );
DFF_X2 U_g1862 ( .D(g1855), .Q(g1862), .CK(CK) );
DFF_X2 U_g1866 ( .D(g1862), .Q(g1866), .CK(CK) );
DFF_X2 U_g1867 ( .D(g24374), .Q(g1867), .CK(CK) );
DFF_X2 U_g1868 ( .D(g24375), .Q(g1868), .CK(CK) );
DFF_X2 U_g1869 ( .D(g24376), .Q(g1869), .CK(CK) );
DFF_X2 U_g1836 ( .D(g25161), .Q(g1836), .CK(CK) );
DFF_X2 U_g1839 ( .D(g25153), .Q(g1839), .CK(CK) );
DFF_X2 U_g1842 ( .D(g25154), .Q(g1842), .CK(CK) );
DFF_X2 U_g1858 ( .D(g25158), .Q(g1858), .CK(CK) );
DFF_X2 U_g1859 ( .D(g25159), .Q(g1859), .CK(CK) );
DFF_X2 U_g1860 ( .D(g25160), .Q(g1860), .CK(CK) );
DFF_X2 U_g1861 ( .D(g24371), .Q(g1861), .CK(CK) );
DFF_X2 U_g1865 ( .D(g24372), .Q(g1865), .CK(CK) );
DFF_X2 U_g1845 ( .D(g24373), .Q(g1845), .CK(CK) );
DFF_X2 U_g1846 ( .D(g25155), .Q(g1846), .CK(CK) );
DFF_X2 U_g1849 ( .D(g25156), .Q(g1849), .CK(CK) );
DFF_X2 U_g1852 ( .D(g25157), .Q(g1852), .CK(CK) );
DFF_X2 U_g1908 ( .D(g16472), .Q(g1908), .CK(CK) );
DFF_X2 U_g1915 ( .D(g1908), .Q(g1915), .CK(CK) );
DFF_X2 U_g1922 ( .D(g1915), .Q(g1922), .CK(CK) );
DFF_X2 U_g1923 ( .D(g19045), .Q(g1923), .CK(CK) );
DFF_X2 U_g1924 ( .D(g1923), .Q(g1924), .CK(CK) );
DFF_X2 U_g1928 ( .D(g29445), .Q(g1928), .CK(CK) );
DFF_X2 U_g1929 ( .D(g19046), .Q(g1929), .CK(CK) );
DFF_X2 U_g1880 ( .D(g1929), .Q(g1880), .CK(CK) );
DFF_X2 U_g1938 ( .D(g19047), .Q(g1938), .CK(CK) );
DFF_X2 U_g1939 ( .D(g1938), .Q(g1939), .CK(CK) );
DFF_X2 U_g1956 ( .D(g28271), .Q(g1956), .CK(CK) );
DFF_X2 U_g1957 ( .D(g28272), .Q(g1957), .CK(CK) );
DFF_X2 U_g1955 ( .D(g28273), .Q(g1955), .CK(CK) );
DFF_X2 U_g1959 ( .D(g28274), .Q(g1959), .CK(CK) );
DFF_X2 U_g1960 ( .D(g28275), .Q(g1960), .CK(CK) );
DFF_X2 U_g1958 ( .D(g28276), .Q(g1958), .CK(CK) );
DFF_X2 U_g1962 ( .D(g28277), .Q(g1962), .CK(CK) );
DFF_X2 U_g1963 ( .D(g28278), .Q(g1963), .CK(CK) );
DFF_X2 U_g1961 ( .D(g28279), .Q(g1961), .CK(CK) );
DFF_X2 U_g1965 ( .D(g28280), .Q(g1965), .CK(CK) );
DFF_X2 U_g1966 ( .D(g28281), .Q(g1966), .CK(CK) );
DFF_X2 U_g1964 ( .D(g28282), .Q(g1964), .CK(CK) );
DFF_X2 U_g1967 ( .D(g26003), .Q(g1967), .CK(CK) );
DFF_X2 U_g1970 ( .D(g26004), .Q(g1970), .CK(CK) );
DFF_X2 U_g1973 ( .D(g26005), .Q(g1973), .CK(CK) );
DFF_X2 U_g1976 ( .D(g26006), .Q(g1976), .CK(CK) );
DFF_X2 U_g1979 ( .D(g26007), .Q(g1979), .CK(CK) );
DFF_X2 U_g1982 ( .D(g26008), .Q(g1982), .CK(CK) );
DFF_X2 U_g1994 ( .D(g29151), .Q(g1994), .CK(CK) );
DFF_X2 U_g1997 ( .D(g29152), .Q(g1997), .CK(CK) );
DFF_X2 U_g2000 ( .D(g29153), .Q(g2000), .CK(CK) );
DFF_X2 U_g1985 ( .D(g29148), .Q(g1985), .CK(CK) );
DFF_X2 U_g1988 ( .D(g29149), .Q(g1988), .CK(CK) );
DFF_X2 U_g1991 ( .D(g29150), .Q(g1991), .CK(CK) );
DFF_X2 U_g1871 ( .D(g27224), .Q(g1871), .CK(CK) );
DFF_X2 U_g1874 ( .D(g27225), .Q(g1874), .CK(CK) );
DFF_X2 U_g1877 ( .D(g27226), .Q(g1877), .CK(CK) );
DFF_X2 U_g1886 ( .D(g8302), .Q(g1886), .CK(CK) );
DFF_X2 U_g1887 ( .D(g24377), .Q(g1887), .CK(CK) );
DFF_X2 U_g1888 ( .D(g19041), .Q(g1888), .CK(CK) );
DFF_X2 U_g1889 ( .D(g19042), .Q(g1889), .CK(CK) );
DFF_X2 U_g1894 ( .D(g19043), .Q(g1894), .CK(CK) );
DFF_X2 U_g1895 ( .D(g19044), .Q(g1895), .CK(CK) );
DFF_X2 U_g1896 ( .D(g29444), .Q(g1896), .CK(CK) );
DFF_X2 U_g1897 ( .D(g29443), .Q(g1897), .CK(CK) );
DFF_X2 U_g1898 ( .D(g29442), .Q(g1898), .CK(CK) );
DFF_X2 U_g1899 ( .D(g29441), .Q(g1899), .CK(CK) );
DFF_X2 U_g1900 ( .D(g29440), .Q(g1900), .CK(CK) );
DFF_X2 U_g1905 ( .D(g1900), .Q(g1905), .CK(CK) );
DFF_X2 U_g1909 ( .D(g13442), .Q(g1909), .CK(CK) );
DFF_X2 U_g1910 ( .D(g13443), .Q(g1910), .CK(CK) );
DFF_X2 U_g1911 ( .D(g13444), .Q(g1911), .CK(CK) );
DFF_X2 U_g1912 ( .D(g13445), .Q(g1912), .CK(CK) );
DFF_X2 U_g1913 ( .D(g13446), .Q(g1913), .CK(CK) );
DFF_X2 U_g1914 ( .D(g13447), .Q(g1914), .CK(CK) );
DFF_X2 U_g1916 ( .D(g13448), .Q(g1916), .CK(CK) );
DFF_X2 U_g1917 ( .D(g13449), .Q(g1917), .CK(CK) );
DFF_X2 U_g1918 ( .D(g26002), .Q(g1918), .CK(CK) );
DFF_X2 U_g1921 ( .D(g13450), .Q(g1921), .CK(CK) );
DFF_X2 U_g2003 ( .D(g13452), .Q(g2003), .CK(CK) );
DFF_X2 U_g2006 ( .D(g2003), .Q(g2006), .CK(CK) );
DFF_X2 U_g2009 ( .D(g2006), .Q(g2009), .CK(CK) );
DFF_X2 U_g2010 ( .D(g20566), .Q(g2010), .CK(CK) );
DFF_X2 U_g2039 ( .D(g21945), .Q(g2039), .CK(CK) );
DFF_X2 U_g2020 ( .D(g23237), .Q(g2020), .CK(CK) );
DFF_X2 U_g2013 ( .D(g24378), .Q(g2013), .CK(CK) );
DFF_X2 U_g2033 ( .D(g25162), .Q(g2033), .CK(CK) );
DFF_X2 U_g2026 ( .D(g26009), .Q(g2026), .CK(CK) );
DFF_X2 U_g2040 ( .D(g26725), .Q(g2040), .CK(CK) );
DFF_X2 U_g2052 ( .D(g27227), .Q(g2052), .CK(CK) );
DFF_X2 U_g2046 ( .D(g27706), .Q(g2046), .CK(CK) );
DFF_X2 U_g2059 ( .D(g28283), .Q(g2059), .CK(CK) );
DFF_X2 U_g2066 ( .D(g28687), .Q(g2066), .CK(CK) );
DFF_X2 U_g2072 ( .D(g29154), .Q(g2072), .CK(CK) );
DFF_X2 U_g2079 ( .D(g23238), .Q(g2079), .CK(CK) );
DFF_X2 U_g2080 ( .D(g23239), .Q(g2080), .CK(CK) );
DFF_X2 U_g2078 ( .D(g23240), .Q(g2078), .CK(CK) );
DFF_X2 U_g2082 ( .D(g23241), .Q(g2082), .CK(CK) );
DFF_X2 U_g2083 ( .D(g23242), .Q(g2083), .CK(CK) );
DFF_X2 U_g2081 ( .D(g23243), .Q(g2081), .CK(CK) );
DFF_X2 U_g2085 ( .D(g23244), .Q(g2085), .CK(CK) );
DFF_X2 U_g2086 ( .D(g23245), .Q(g2086), .CK(CK) );
DFF_X2 U_g2084 ( .D(g23246), .Q(g2084), .CK(CK) );
DFF_X2 U_g2088 ( .D(g23247), .Q(g2088), .CK(CK) );
DFF_X2 U_g2089 ( .D(g23248), .Q(g2089), .CK(CK) );
DFF_X2 U_g2087 ( .D(g23249), .Q(g2087), .CK(CK) );
DFF_X2 U_g2091 ( .D(g23250), .Q(g2091), .CK(CK) );
DFF_X2 U_g2092 ( .D(g23251), .Q(g2092), .CK(CK) );
DFF_X2 U_g2090 ( .D(g23252), .Q(g2090), .CK(CK) );
DFF_X2 U_g2094 ( .D(g23253), .Q(g2094), .CK(CK) );
DFF_X2 U_g2095 ( .D(g23254), .Q(g2095), .CK(CK) );
DFF_X2 U_g2093 ( .D(g23255), .Q(g2093), .CK(CK) );
DFF_X2 U_g2097 ( .D(g23256), .Q(g2097), .CK(CK) );
DFF_X2 U_g2098 ( .D(g23257), .Q(g2098), .CK(CK) );
DFF_X2 U_g2096 ( .D(g23258), .Q(g2096), .CK(CK) );
DFF_X2 U_g2100 ( .D(g23259), .Q(g2100), .CK(CK) );
DFF_X2 U_g2101 ( .D(g23260), .Q(g2101), .CK(CK) );
DFF_X2 U_g2099 ( .D(g23261), .Q(g2099), .CK(CK) );
DFF_X2 U_g2103 ( .D(g23262), .Q(g2103), .CK(CK) );
DFF_X2 U_g2104 ( .D(g23263), .Q(g2104), .CK(CK) );
DFF_X2 U_g2102 ( .D(g23264), .Q(g2102), .CK(CK) );
DFF_X2 U_g2106 ( .D(g23265), .Q(g2106), .CK(CK) );
DFF_X2 U_g2107 ( .D(g23266), .Q(g2107), .CK(CK) );
DFF_X2 U_g2105 ( .D(g23267), .Q(g2105), .CK(CK) );
DFF_X2 U_g2109 ( .D(g23268), .Q(g2109), .CK(CK) );
DFF_X2 U_g2110 ( .D(g23269), .Q(g2110), .CK(CK) );
DFF_X2 U_g2108 ( .D(g23270), .Q(g2108), .CK(CK) );
DFF_X2 U_g2112 ( .D(g23271), .Q(g2112), .CK(CK) );
DFF_X2 U_g2113 ( .D(g23272), .Q(g2113), .CK(CK) );
DFF_X2 U_g2111 ( .D(g23273), .Q(g2111), .CK(CK) );
DFF_X2 U_g2115 ( .D(g26726), .Q(g2115), .CK(CK) );
DFF_X2 U_g2116 ( .D(g26727), .Q(g2116), .CK(CK) );
DFF_X2 U_g2114 ( .D(g26728), .Q(g2114), .CK(CK) );
DFF_X2 U_g2118 ( .D(g24379), .Q(g2118), .CK(CK) );
DFF_X2 U_g2119 ( .D(g24380), .Q(g2119), .CK(CK) );
DFF_X2 U_g2117 ( .D(g24381), .Q(g2117), .CK(CK) );
DFF_X2 U_g2214 ( .D(g13453), .Q(g2214), .CK(CK) );
DFF_X2 U_g2211 ( .D(g2214), .Q(g2211), .CK(CK) );
DFF_X2 U_g2241 ( .D(g2211), .Q(g2241), .CK(CK) );
DFF_X2 U_g2206 ( .D(g24382), .Q(g2206), .CK(CK) );
DFF_X2 U_g2207 ( .D(g24383), .Q(g2207), .CK(CK) );
DFF_X2 U_g2205 ( .D(g24384), .Q(g2205), .CK(CK) );
DFF_X2 U_g2209 ( .D(g24385), .Q(g2209), .CK(CK) );
DFF_X2 U_g2210 ( .D(g24386), .Q(g2210), .CK(CK) );
DFF_X2 U_g2208 ( .D(g24387), .Q(g2208), .CK(CK) );
DFF_X2 U_g2218 ( .D(g24388), .Q(g2218), .CK(CK) );
DFF_X2 U_g2219 ( .D(g24389), .Q(g2219), .CK(CK) );
DFF_X2 U_g2217 ( .D(g24390), .Q(g2217), .CK(CK) );
DFF_X2 U_g2221 ( .D(g24391), .Q(g2221), .CK(CK) );
DFF_X2 U_g2222 ( .D(g24392), .Q(g2222), .CK(CK) );
DFF_X2 U_g2220 ( .D(g24393), .Q(g2220), .CK(CK) );
DFF_X2 U_g2224 ( .D(g24394), .Q(g2224), .CK(CK) );
DFF_X2 U_g2225 ( .D(g24395), .Q(g2225), .CK(CK) );
DFF_X2 U_g2223 ( .D(g24396), .Q(g2223), .CK(CK) );
DFF_X2 U_g2227 ( .D(g24397), .Q(g2227), .CK(CK) );
DFF_X2 U_g2228 ( .D(g24398), .Q(g2228), .CK(CK) );
DFF_X2 U_g2226 ( .D(g24399), .Q(g2226), .CK(CK) );
DFF_X2 U_g2230 ( .D(g24400), .Q(g2230), .CK(CK) );
DFF_X2 U_g2231 ( .D(g24401), .Q(g2231), .CK(CK) );
DFF_X2 U_g2229 ( .D(g24402), .Q(g2229), .CK(CK) );
DFF_X2 U_g2233 ( .D(g24403), .Q(g2233), .CK(CK) );
DFF_X2 U_g2234 ( .D(g24404), .Q(g2234), .CK(CK) );
DFF_X2 U_g2232 ( .D(g24405), .Q(g2232), .CK(CK) );
DFF_X2 U_g2236 ( .D(g24406), .Q(g2236), .CK(CK) );
DFF_X2 U_g2237 ( .D(g24407), .Q(g2237), .CK(CK) );
DFF_X2 U_g2235 ( .D(g24408), .Q(g2235), .CK(CK) );
DFF_X2 U_g2239 ( .D(g24409), .Q(g2239), .CK(CK) );
DFF_X2 U_g2240 ( .D(g24410), .Q(g2240), .CK(CK) );
DFF_X2 U_g2238 ( .D(g24411), .Q(g2238), .CK(CK) );
DFF_X2 U_g2245 ( .D(g26730), .Q(g2245), .CK(CK) );
DFF_X2 U_g2246 ( .D(g26731), .Q(g2246), .CK(CK) );
DFF_X2 U_g2244 ( .D(g26732), .Q(g2244), .CK(CK) );
DFF_X2 U_g2248 ( .D(g26733), .Q(g2248), .CK(CK) );
DFF_X2 U_g2249 ( .D(g26734), .Q(g2249), .CK(CK) );
DFF_X2 U_g2247 ( .D(g26735), .Q(g2247), .CK(CK) );
DFF_X2 U_g2251 ( .D(g26736), .Q(g2251), .CK(CK) );
DFF_X2 U_g2252 ( .D(g26737), .Q(g2252), .CK(CK) );
DFF_X2 U_g2250 ( .D(g26738), .Q(g2250), .CK(CK) );
DFF_X2 U_g2254 ( .D(g26739), .Q(g2254), .CK(CK) );
DFF_X2 U_g2255 ( .D(g26740), .Q(g2255), .CK(CK) );
DFF_X2 U_g2253 ( .D(g26741), .Q(g2253), .CK(CK) );
DFF_X2 U_g2261 ( .D(g30551), .Q(g2261), .CK(CK) );
DFF_X2 U_g2264 ( .D(g30552), .Q(g2264), .CK(CK) );
DFF_X2 U_g2267 ( .D(g30553), .Q(g2267), .CK(CK) );
DFF_X2 U_g2306 ( .D(g30896), .Q(g2306), .CK(CK) );
DFF_X2 U_g2309 ( .D(g30897), .Q(g2309), .CK(CK) );
DFF_X2 U_g2312 ( .D(g30898), .Q(g2312), .CK(CK) );
DFF_X2 U_g2270 ( .D(g30890), .Q(g2270), .CK(CK) );
DFF_X2 U_g2273 ( .D(g30891), .Q(g2273), .CK(CK) );
DFF_X2 U_g2276 ( .D(g30892), .Q(g2276), .CK(CK) );
DFF_X2 U_g2315 ( .D(g30899), .Q(g2315), .CK(CK) );
DFF_X2 U_g2318 ( .D(g30900), .Q(g2318), .CK(CK) );
DFF_X2 U_g2321 ( .D(g30901), .Q(g2321), .CK(CK) );
DFF_X2 U_g2279 ( .D(g30554), .Q(g2279), .CK(CK) );
DFF_X2 U_g2282 ( .D(g30555), .Q(g2282), .CK(CK) );
DFF_X2 U_g2285 ( .D(g30556), .Q(g2285), .CK(CK) );
DFF_X2 U_g2324 ( .D(g30560), .Q(g2324), .CK(CK) );
DFF_X2 U_g2327 ( .D(g30561), .Q(g2327), .CK(CK) );
DFF_X2 U_g2330 ( .D(g30562), .Q(g2330), .CK(CK) );
DFF_X2 U_g2288 ( .D(g30557), .Q(g2288), .CK(CK) );
DFF_X2 U_g2291 ( .D(g30558), .Q(g2291), .CK(CK) );
DFF_X2 U_g2294 ( .D(g30559), .Q(g2294), .CK(CK) );
DFF_X2 U_g2333 ( .D(g30563), .Q(g2333), .CK(CK) );
DFF_X2 U_g2336 ( .D(g30564), .Q(g2336), .CK(CK) );
DFF_X2 U_g2339 ( .D(g30565), .Q(g2339), .CK(CK) );
DFF_X2 U_g2297 ( .D(g30893), .Q(g2297), .CK(CK) );
DFF_X2 U_g2300 ( .D(g30894), .Q(g2300), .CK(CK) );
DFF_X2 U_g2303 ( .D(g30895), .Q(g2303), .CK(CK) );
DFF_X2 U_g2342 ( .D(g30902), .Q(g2342), .CK(CK) );
DFF_X2 U_g2345 ( .D(g30903), .Q(g2345), .CK(CK) );
DFF_X2 U_g2348 ( .D(g30904), .Q(g2348), .CK(CK) );
DFF_X2 U_g2160 ( .D(g26010), .Q(g2160), .CK(CK) );
DFF_X2 U_g2156 ( .D(g26729), .Q(g2156), .CK(CK) );
DFF_X2 U_g2151 ( .D(g27228), .Q(g2151), .CK(CK) );
DFF_X2 U_g2147 ( .D(g27707), .Q(g2147), .CK(CK) );
DFF_X2 U_g2142 ( .D(g28284), .Q(g2142), .CK(CK) );
DFF_X2 U_g2138 ( .D(g28688), .Q(g2138), .CK(CK) );
DFF_X2 U_g2133 ( .D(g29155), .Q(g2133), .CK(CK) );
DFF_X2 U_g2129 ( .D(g29446), .Q(g2129), .CK(CK) );
DFF_X2 U_g2124 ( .D(g29648), .Q(g2124), .CK(CK) );
DFF_X2 U_g2120 ( .D(g29806), .Q(g2120), .CK(CK) );
DFF_X2 U_g2256 ( .D(g20567), .Q(g2256), .CK(CK) );
DFF_X2 U_g2258 ( .D(g2256), .Q(g2258), .CK(CK) );
DFF_X2 U_g2257 ( .D(g2258), .Q(g2257), .CK(CK) );
DFF_X2 U_g2351 ( .D(g13454), .Q(g2351), .CK(CK) );
DFF_X2 U_g2480 ( .D(g2351), .Q(g2480), .CK(CK) );
DFF_X2 U_g2476 ( .D(g2480), .Q(g2476), .CK(CK) );
DFF_X2 U_g2384 ( .D(g11577), .Q(g2384), .CK(CK) );
DFF_X2 U_g2429 ( .D(g28285), .Q(g2429), .CK(CK) );
DFF_X2 U_g2418 ( .D(g28286), .Q(g2418), .CK(CK) );
DFF_X2 U_g2421 ( .D(g28287), .Q(g2421), .CK(CK) );
DFF_X2 U_g2444 ( .D(g28288), .Q(g2444), .CK(CK) );
DFF_X2 U_g2433 ( .D(g28289), .Q(g2433), .CK(CK) );
DFF_X2 U_g2436 ( .D(g28290), .Q(g2436), .CK(CK) );
DFF_X2 U_g2459 ( .D(g28291), .Q(g2459), .CK(CK) );
DFF_X2 U_g2448 ( .D(g28292), .Q(g2448), .CK(CK) );
DFF_X2 U_g2451 ( .D(g28293), .Q(g2451), .CK(CK) );
DFF_X2 U_g2473 ( .D(g28294), .Q(g2473), .CK(CK) );
DFF_X2 U_g2463 ( .D(g28295), .Q(g2463), .CK(CK) );
DFF_X2 U_g2466 ( .D(g28296), .Q(g2466), .CK(CK) );
DFF_X2 U_g2483 ( .D(g29447), .Q(g2483), .CK(CK) );
DFF_X2 U_g2486 ( .D(g29448), .Q(g2486), .CK(CK) );
DFF_X2 U_g2489 ( .D(g29449), .Q(g2489), .CK(CK) );
DFF_X2 U_g2492 ( .D(g29652), .Q(g2492), .CK(CK) );
DFF_X2 U_g2495 ( .D(g29653), .Q(g2495), .CK(CK) );
DFF_X2 U_g2498 ( .D(g29654), .Q(g2498), .CK(CK) );
DFF_X2 U_g2502 ( .D(g29450), .Q(g2502), .CK(CK) );
DFF_X2 U_g2503 ( .D(g29451), .Q(g2503), .CK(CK) );
DFF_X2 U_g2501 ( .D(g29452), .Q(g2501), .CK(CK) );
DFF_X2 U_g2504 ( .D(g27708), .Q(g2504), .CK(CK) );
DFF_X2 U_g2507 ( .D(g27709), .Q(g2507), .CK(CK) );
DFF_X2 U_g2510 ( .D(g27710), .Q(g2510), .CK(CK) );
DFF_X2 U_g2513 ( .D(g27711), .Q(g2513), .CK(CK) );
DFF_X2 U_g2516 ( .D(g27712), .Q(g2516), .CK(CK) );
DFF_X2 U_g2519 ( .D(g27713), .Q(g2519), .CK(CK) );
DFF_X2 U_g2523 ( .D(g28689), .Q(g2523), .CK(CK) );
DFF_X2 U_g2524 ( .D(g28690), .Q(g2524), .CK(CK) );
DFF_X2 U_g2522 ( .D(g28691), .Q(g2522), .CK(CK) );
DFF_X2 U_g2387 ( .D(g29807), .Q(g2387), .CK(CK) );
DFF_X2 U_g2388 ( .D(g29808), .Q(g2388), .CK(CK) );
DFF_X2 U_g2389 ( .D(g29809), .Q(g2389), .CK(CK) );
DFF_X2 U_g2390 ( .D(g30905), .Q(g2390), .CK(CK) );
DFF_X2 U_g2391 ( .D(g30906), .Q(g2391), .CK(CK) );
DFF_X2 U_g2392 ( .D(g30907), .Q(g2392), .CK(CK) );
DFF_X2 U_g2393 ( .D(g30719), .Q(g2393), .CK(CK) );
DFF_X2 U_g2394 ( .D(g30720), .Q(g2394), .CK(CK) );
DFF_X2 U_g2395 ( .D(g30721), .Q(g2395), .CK(CK) );
DFF_X2 U_g2397 ( .D(g29649), .Q(g2397), .CK(CK) );
DFF_X2 U_g2398 ( .D(g29650), .Q(g2398), .CK(CK) );
DFF_X2 U_g2396 ( .D(g29651), .Q(g2396), .CK(CK) );
DFF_X2 U_g2478 ( .D(g27230), .Q(g2478), .CK(CK) );
DFF_X2 U_g2479 ( .D(g27231), .Q(g2479), .CK(CK) );
DFF_X2 U_g2477 ( .D(g27232), .Q(g2477), .CK(CK) );
DFF_X2 U_g2525 ( .D(g11590), .Q(g2525), .CK(CK) );
DFF_X2 U_g2526 ( .D(g2525), .Q(g2526), .CK(CK) );
DFF_X2 U_g2527 ( .D(g11591), .Q(g2527), .CK(CK) );
DFF_X2 U_g2528 ( .D(g2527), .Q(g2528), .CK(CK) );
DFF_X2 U_g2529 ( .D(g11592), .Q(g2529), .CK(CK) );
DFF_X2 U_g2354 ( .D(g2529), .Q(g2354), .CK(CK) );
DFF_X2 U_g2355 ( .D(g11572), .Q(g2355), .CK(CK) );
DFF_X2 U_g2356 ( .D(g2355), .Q(g2356), .CK(CK) );
DFF_X2 U_g2357 ( .D(g11573), .Q(g2357), .CK(CK) );
DFF_X2 U_g2358 ( .D(g2357), .Q(g2358), .CK(CK) );
DFF_X2 U_g2359 ( .D(g11574), .Q(g2359), .CK(CK) );
DFF_X2 U_g2360 ( .D(g2359), .Q(g2360), .CK(CK) );
DFF_X2 U_g2361 ( .D(g11575), .Q(g2361), .CK(CK) );
DFF_X2 U_g2362 ( .D(g2361), .Q(g2362), .CK(CK) );
DFF_X2 U_g2363 ( .D(g11576), .Q(g2363), .CK(CK) );
DFF_X2 U_g2364 ( .D(g2363), .Q(g2364), .CK(CK) );
DFF_X2 U_g2365 ( .D(g13455), .Q(g2365), .CK(CK) );
DFF_X2 U_g2366 ( .D(g2365), .Q(g2366), .CK(CK) );
DFF_X2 U_g2374 ( .D(g19048), .Q(g2374), .CK(CK) );
DFF_X2 U_g2380 ( .D(g30314), .Q(g2380), .CK(CK) );
DFF_X2 U_g2383 ( .D(g30315), .Q(g2383), .CK(CK) );
DFF_X2 U_g2372 ( .D(g30316), .Q(g2372), .CK(CK) );
DFF_X2 U_g2371 ( .D(g30317), .Q(g2371), .CK(CK) );
DFF_X2 U_g2370 ( .D(g30318), .Q(g2370), .CK(CK) );
DFF_X2 U_g2369 ( .D(g30319), .Q(g2369), .CK(CK) );
DFF_X2 U_g2379 ( .D(g19052), .Q(g2379), .CK(CK) );
DFF_X2 U_g2378 ( .D(g19051), .Q(g2378), .CK(CK) );
DFF_X2 U_g2377 ( .D(g19050), .Q(g2377), .CK(CK) );
DFF_X2 U_g2376 ( .D(g19049), .Q(g2376), .CK(CK) );
DFF_X2 U_g2375 ( .D(g25163), .Q(g2375), .CK(CK) );
DFF_X2 U_g2373 ( .D(g27229), .Q(g2373), .CK(CK) );
DFF_X2 U_g2417 ( .D(g11578), .Q(g2417), .CK(CK) );
DFF_X2 U_g2424 ( .D(g2417), .Q(g2424), .CK(CK) );
DFF_X2 U_g2425 ( .D(g11579), .Q(g2425), .CK(CK) );
DFF_X2 U_g2426 ( .D(g2425), .Q(g2426), .CK(CK) );
DFF_X2 U_g2427 ( .D(g11580), .Q(g2427), .CK(CK) );
DFF_X2 U_g2428 ( .D(g2427), .Q(g2428), .CK(CK) );
DFF_X2 U_g2432 ( .D(g11581), .Q(g2432), .CK(CK) );
DFF_X2 U_g2439 ( .D(g2432), .Q(g2439), .CK(CK) );
DFF_X2 U_g2440 ( .D(g11582), .Q(g2440), .CK(CK) );
DFF_X2 U_g2441 ( .D(g2440), .Q(g2441), .CK(CK) );
DFF_X2 U_g2442 ( .D(g11583), .Q(g2442), .CK(CK) );
DFF_X2 U_g2443 ( .D(g2442), .Q(g2443), .CK(CK) );
DFF_X2 U_g2447 ( .D(g11584), .Q(g2447), .CK(CK) );
DFF_X2 U_g2454 ( .D(g2447), .Q(g2454), .CK(CK) );
DFF_X2 U_g2455 ( .D(g11585), .Q(g2455), .CK(CK) );
DFF_X2 U_g2456 ( .D(g2455), .Q(g2456), .CK(CK) );
DFF_X2 U_g2457 ( .D(g11586), .Q(g2457), .CK(CK) );
DFF_X2 U_g2458 ( .D(g2457), .Q(g2458), .CK(CK) );
DFF_X2 U_g2462 ( .D(g11587), .Q(g2462), .CK(CK) );
DFF_X2 U_g2469 ( .D(g2462), .Q(g2469), .CK(CK) );
DFF_X2 U_g2470 ( .D(g11588), .Q(g2470), .CK(CK) );
DFF_X2 U_g2471 ( .D(g2470), .Q(g2471), .CK(CK) );
DFF_X2 U_g2472 ( .D(g11589), .Q(g2472), .CK(CK) );
DFF_X2 U_g2399 ( .D(g2472), .Q(g2399), .CK(CK) );
DFF_X2 U_g2400 ( .D(g13456), .Q(g2400), .CK(CK) );
DFF_X2 U_g2406 ( .D(g2400), .Q(g2406), .CK(CK) );
DFF_X2 U_g2412 ( .D(g2406), .Q(g2412), .CK(CK) );
DFF_X2 U_g2619 ( .D(g13467), .Q(g2619), .CK(CK) );
DFF_X2 U_g2625 ( .D(g2619), .Q(g2625), .CK(CK) );
DFF_X2 U_g2624 ( .D(g2625), .Q(g2624), .CK(CK) );
DFF_X2 U_g2628 ( .D(g23274), .Q(g2628), .CK(CK) );
DFF_X2 U_g2631 ( .D(g20568), .Q(g2631), .CK(CK) );
DFF_X2 U_g2584 ( .D(g20569), .Q(g2584), .CK(CK) );
DFF_X2 U_g2587 ( .D(g16473), .Q(g2587), .CK(CK) );
DFF_X2 U_g2597 ( .D(g2587), .Q(g2597), .CK(CK) );
DFF_X2 U_g2598 ( .D(g2597), .Q(g2598), .CK(CK) );
DFF_X2 U_g2638 ( .D(g11593), .Q(g2638), .CK(CK) );
DFF_X2 U_g2643 ( .D(g2638), .Q(g2643), .CK(CK) );
DFF_X2 U_g2644 ( .D(g11596), .Q(g2644), .CK(CK) );
DFF_X2 U_g2645 ( .D(g2644), .Q(g2645), .CK(CK) );
DFF_X2 U_g2646 ( .D(g11597), .Q(g2646), .CK(CK) );
DFF_X2 U_g2647 ( .D(g2646), .Q(g2647), .CK(CK) );
DFF_X2 U_g2648 ( .D(g11598), .Q(g2648), .CK(CK) );
DFF_X2 U_g2639 ( .D(g2648), .Q(g2639), .CK(CK) );
DFF_X2 U_g2640 ( .D(g11594), .Q(g2640), .CK(CK) );
DFF_X2 U_g2641 ( .D(g2640), .Q(g2641), .CK(CK) );
DFF_X2 U_g2642 ( .D(g11595), .Q(g2642), .CK(CK) );
DFF_X2 U_g2564 ( .D(g2642), .Q(g2564), .CK(CK) );
DFF_X2 U_g2549 ( .D(g13457), .Q(g2549), .CK(CK) );
DFF_X2 U_g2556 ( .D(g2549), .Q(g2556), .CK(CK) );
DFF_X2 U_g2560 ( .D(g2556), .Q(g2560), .CK(CK) );
DFF_X2 U_g2561 ( .D(g24415), .Q(g2561), .CK(CK) );
DFF_X2 U_g2562 ( .D(g24416), .Q(g2562), .CK(CK) );
DFF_X2 U_g2563 ( .D(g24417), .Q(g2563), .CK(CK) );
DFF_X2 U_g2530 ( .D(g25172), .Q(g2530), .CK(CK) );
DFF_X2 U_g2533 ( .D(g25164), .Q(g2533), .CK(CK) );
DFF_X2 U_g2536 ( .D(g25165), .Q(g2536), .CK(CK) );
DFF_X2 U_g2552 ( .D(g25169), .Q(g2552), .CK(CK) );
DFF_X2 U_g2553 ( .D(g25170), .Q(g2553), .CK(CK) );
DFF_X2 U_g2554 ( .D(g25171), .Q(g2554), .CK(CK) );
DFF_X2 U_g2555 ( .D(g24412), .Q(g2555), .CK(CK) );
DFF_X2 U_g2559 ( .D(g24413), .Q(g2559), .CK(CK) );
DFF_X2 U_g2539 ( .D(g24414), .Q(g2539), .CK(CK) );
DFF_X2 U_g2540 ( .D(g25166), .Q(g2540), .CK(CK) );
DFF_X2 U_g2543 ( .D(g25167), .Q(g2543), .CK(CK) );
DFF_X2 U_g2546 ( .D(g25168), .Q(g2546), .CK(CK) );
DFF_X2 U_g2602 ( .D(g16474), .Q(g2602), .CK(CK) );
DFF_X2 U_g2609 ( .D(g2602), .Q(g2609), .CK(CK) );
DFF_X2 U_g2616 ( .D(g2609), .Q(g2616), .CK(CK) );
DFF_X2 U_g2617 ( .D(g19057), .Q(g2617), .CK(CK) );
DFF_X2 U_g2618 ( .D(g2617), .Q(g2618), .CK(CK) );
DFF_X2 U_g2622 ( .D(g30325), .Q(g2622), .CK(CK) );
DFF_X2 U_g2623 ( .D(g19058), .Q(g2623), .CK(CK) );
DFF_X2 U_g2574 ( .D(g2623), .Q(g2574), .CK(CK) );
DFF_X2 U_g2632 ( .D(g19059), .Q(g2632), .CK(CK) );
DFF_X2 U_g2633 ( .D(g2632), .Q(g2633), .CK(CK) );
DFF_X2 U_g2650 ( .D(g28297), .Q(g2650), .CK(CK) );
DFF_X2 U_g2651 ( .D(g28298), .Q(g2651), .CK(CK) );
DFF_X2 U_g2649 ( .D(g28299), .Q(g2649), .CK(CK) );
DFF_X2 U_g2653 ( .D(g28300), .Q(g2653), .CK(CK) );
DFF_X2 U_g2654 ( .D(g28301), .Q(g2654), .CK(CK) );
DFF_X2 U_g2652 ( .D(g28302), .Q(g2652), .CK(CK) );
DFF_X2 U_g2656 ( .D(g28303), .Q(g2656), .CK(CK) );
DFF_X2 U_g2657 ( .D(g28304), .Q(g2657), .CK(CK) );
DFF_X2 U_g2655 ( .D(g28305), .Q(g2655), .CK(CK) );
DFF_X2 U_g2659 ( .D(g28306), .Q(g2659), .CK(CK) );
DFF_X2 U_g2660 ( .D(g28307), .Q(g2660), .CK(CK) );
DFF_X2 U_g2658 ( .D(g28308), .Q(g2658), .CK(CK) );
DFF_X2 U_g2661 ( .D(g26012), .Q(g2661), .CK(CK) );
DFF_X2 U_g2664 ( .D(g26013), .Q(g2664), .CK(CK) );
DFF_X2 U_g2667 ( .D(g26014), .Q(g2667), .CK(CK) );
DFF_X2 U_g2670 ( .D(g26015), .Q(g2670), .CK(CK) );
DFF_X2 U_g2673 ( .D(g26016), .Q(g2673), .CK(CK) );
DFF_X2 U_g2676 ( .D(g26017), .Q(g2676), .CK(CK) );
DFF_X2 U_g2688 ( .D(g29159), .Q(g2688), .CK(CK) );
DFF_X2 U_g2691 ( .D(g29160), .Q(g2691), .CK(CK) );
DFF_X2 U_g2694 ( .D(g29161), .Q(g2694), .CK(CK) );
DFF_X2 U_g2679 ( .D(g29156), .Q(g2679), .CK(CK) );
DFF_X2 U_g2682 ( .D(g29157), .Q(g2682), .CK(CK) );
DFF_X2 U_g2685 ( .D(g29158), .Q(g2685), .CK(CK) );
DFF_X2 U_g2565 ( .D(g27233), .Q(g2565), .CK(CK) );
DFF_X2 U_g2568 ( .D(g27234), .Q(g2568), .CK(CK) );
DFF_X2 U_g2571 ( .D(g27235), .Q(g2571), .CK(CK) );
DFF_X2 U_g2580 ( .D(g8311), .Q(g2580), .CK(CK) );
DFF_X2 U_g2581 ( .D(g24418), .Q(g2581), .CK(CK) );
DFF_X2 U_g2582 ( .D(g19053), .Q(g2582), .CK(CK) );
DFF_X2 U_g2583 ( .D(g19054), .Q(g2583), .CK(CK) );
DFF_X2 U_g2588 ( .D(g19055), .Q(g2588), .CK(CK) );
DFF_X2 U_g2589 ( .D(g19056), .Q(g2589), .CK(CK) );
DFF_X2 U_g2590 ( .D(g30324), .Q(g2590), .CK(CK) );
DFF_X2 U_g2591 ( .D(g30323), .Q(g2591), .CK(CK) );
DFF_X2 U_g2592 ( .D(g30322), .Q(g2592), .CK(CK) );
DFF_X2 U_g2593 ( .D(g30321), .Q(g2593), .CK(CK) );
DFF_X2 U_g2594 ( .D(g30320), .Q(g2594), .CK(CK) );
DFF_X2 U_g2599 ( .D(g2594), .Q(g2599), .CK(CK) );
DFF_X2 U_g2603 ( .D(g13458), .Q(g2603), .CK(CK) );
DFF_X2 U_g2604 ( .D(g13459), .Q(g2604), .CK(CK) );
DFF_X2 U_g2605 ( .D(g13460), .Q(g2605), .CK(CK) );
DFF_X2 U_g2606 ( .D(g13461), .Q(g2606), .CK(CK) );
DFF_X2 U_g2607 ( .D(g13462), .Q(g2607), .CK(CK) );
DFF_X2 U_g2608 ( .D(g13463), .Q(g2608), .CK(CK) );
DFF_X2 U_g2610 ( .D(g13464), .Q(g2610), .CK(CK) );
DFF_X2 U_g2611 ( .D(g13465), .Q(g2611), .CK(CK) );
DFF_X2 U_g2612 ( .D(g26011), .Q(g2612), .CK(CK) );
DFF_X2 U_g2615 ( .D(g13466), .Q(g2615), .CK(CK) );
DFF_X2 U_g2697 ( .D(g13468), .Q(g2697), .CK(CK) );
DFF_X2 U_g2700 ( .D(g2697), .Q(g2700), .CK(CK) );
DFF_X2 U_g2703 ( .D(g2700), .Q(g2703), .CK(CK) );
DFF_X2 U_g2704 ( .D(g20570), .Q(g2704), .CK(CK) );
DFF_X2 U_g2733 ( .D(g21946), .Q(g2733), .CK(CK) );
DFF_X2 U_g2714 ( .D(g23275), .Q(g2714), .CK(CK) );
DFF_X2 U_g2707 ( .D(g24419), .Q(g2707), .CK(CK) );
DFF_X2 U_g2727 ( .D(g25173), .Q(g2727), .CK(CK) );
DFF_X2 U_g2720 ( .D(g26018), .Q(g2720), .CK(CK) );
DFF_X2 U_g2734 ( .D(g26742), .Q(g2734), .CK(CK) );
DFF_X2 U_g2746 ( .D(g27236), .Q(g2746), .CK(CK) );
DFF_X2 U_g2740 ( .D(g27714), .Q(g2740), .CK(CK) );
DFF_X2 U_g2753 ( .D(g28309), .Q(g2753), .CK(CK) );
DFF_X2 U_g2760 ( .D(g28692), .Q(g2760), .CK(CK) );
DFF_X2 U_g2766 ( .D(g29162), .Q(g2766), .CK(CK) );
DFF_X2 U_g2773 ( .D(g23276), .Q(g2773), .CK(CK) );
DFF_X2 U_g2774 ( .D(g23277), .Q(g2774), .CK(CK) );
DFF_X2 U_g2772 ( .D(g23278), .Q(g2772), .CK(CK) );
DFF_X2 U_g2776 ( .D(g23279), .Q(g2776), .CK(CK) );
DFF_X2 U_g2777 ( .D(g23280), .Q(g2777), .CK(CK) );
DFF_X2 U_g2775 ( .D(g23281), .Q(g2775), .CK(CK) );
DFF_X2 U_g2779 ( .D(g23282), .Q(g2779), .CK(CK) );
DFF_X2 U_g2780 ( .D(g23283), .Q(g2780), .CK(CK) );
DFF_X2 U_g2778 ( .D(g23284), .Q(g2778), .CK(CK) );
DFF_X2 U_g2782 ( .D(g23285), .Q(g2782), .CK(CK) );
DFF_X2 U_g2783 ( .D(g23286), .Q(g2783), .CK(CK) );
DFF_X2 U_g2781 ( .D(g23287), .Q(g2781), .CK(CK) );
DFF_X2 U_g2785 ( .D(g23288), .Q(g2785), .CK(CK) );
DFF_X2 U_g2786 ( .D(g23289), .Q(g2786), .CK(CK) );
DFF_X2 U_g2784 ( .D(g23290), .Q(g2784), .CK(CK) );
DFF_X2 U_g2788 ( .D(g23291), .Q(g2788), .CK(CK) );
DFF_X2 U_g2789 ( .D(g23292), .Q(g2789), .CK(CK) );
DFF_X2 U_g2787 ( .D(g23293), .Q(g2787), .CK(CK) );
DFF_X2 U_g2791 ( .D(g23294), .Q(g2791), .CK(CK) );
DFF_X2 U_g2792 ( .D(g23295), .Q(g2792), .CK(CK) );
DFF_X2 U_g2790 ( .D(g23296), .Q(g2790), .CK(CK) );
DFF_X2 U_g2794 ( .D(g23297), .Q(g2794), .CK(CK) );
DFF_X2 U_g2795 ( .D(g23298), .Q(g2795), .CK(CK) );
DFF_X2 U_g2793 ( .D(g23299), .Q(g2793), .CK(CK) );
DFF_X2 U_g2797 ( .D(g23300), .Q(g2797), .CK(CK) );
DFF_X2 U_g2798 ( .D(g23301), .Q(g2798), .CK(CK) );
DFF_X2 U_g2796 ( .D(g23302), .Q(g2796), .CK(CK) );
DFF_X2 U_g2800 ( .D(g23303), .Q(g2800), .CK(CK) );
DFF_X2 U_g2801 ( .D(g23304), .Q(g2801), .CK(CK) );
DFF_X2 U_g2799 ( .D(g23305), .Q(g2799), .CK(CK) );
DFF_X2 U_g2803 ( .D(g23306), .Q(g2803), .CK(CK) );
DFF_X2 U_g2804 ( .D(g23307), .Q(g2804), .CK(CK) );
DFF_X2 U_g2802 ( .D(g23308), .Q(g2802), .CK(CK) );
DFF_X2 U_g2806 ( .D(g23309), .Q(g2806), .CK(CK) );
DFF_X2 U_g2807 ( .D(g23310), .Q(g2807), .CK(CK) );
DFF_X2 U_g2805 ( .D(g23311), .Q(g2805), .CK(CK) );
DFF_X2 U_g2809 ( .D(g26743), .Q(g2809), .CK(CK) );
DFF_X2 U_g2810 ( .D(g26744), .Q(g2810), .CK(CK) );
DFF_X2 U_g2808 ( .D(g26745), .Q(g2808), .CK(CK) );
DFF_X2 U_g2812 ( .D(g24420), .Q(g2812), .CK(CK) );
DFF_X2 U_g2813 ( .D(g24421), .Q(g2813), .CK(CK) );
DFF_X2 U_g2811 ( .D(g24422), .Q(g2811), .CK(CK) );
DFF_X2 U_g3054 ( .D(g23317), .Q(g3054), .CK(CK) );
DFF_X2 U_g3079 ( .D(g23318), .Q(g3079), .CK(CK) );
DFF_X2 U_g3080 ( .D(g21965), .Q(g3080), .CK(CK) );
DFF_X2 U_g3043 ( .D(g29453), .Q(g3043), .CK(CK) );
DFF_X2 U_g3044 ( .D(g29454), .Q(g3044), .CK(CK) );
DFF_X2 U_g3045 ( .D(g29455), .Q(g3045), .CK(CK) );
DFF_X2 U_g3046 ( .D(g29456), .Q(g3046), .CK(CK) );
DFF_X2 U_g3047 ( .D(g29457), .Q(g3047), .CK(CK) );
DFF_X2 U_g3048 ( .D(g29458), .Q(g3048), .CK(CK) );
DFF_X2 U_g3049 ( .D(g29459), .Q(g3049), .CK(CK) );
DFF_X2 U_g3050 ( .D(g29460), .Q(g3050), .CK(CK) );
DFF_X2 U_g3051 ( .D(g29655), .Q(g3051), .CK(CK) );
DFF_X2 U_g3052 ( .D(g29972), .Q(g3052), .CK(CK) );
DFF_X2 U_g3053 ( .D(g29973), .Q(g3053), .CK(CK) );
DFF_X2 U_g3055 ( .D(g29974), .Q(g3055), .CK(CK) );
DFF_X2 U_g3056 ( .D(g29975), .Q(g3056), .CK(CK) );
DFF_X2 U_g3057 ( .D(g29976), .Q(g3057), .CK(CK) );
DFF_X2 U_g3058 ( .D(g29977), .Q(g3058), .CK(CK) );
DFF_X2 U_g3059 ( .D(g29978), .Q(g3059), .CK(CK) );
DFF_X2 U_g3060 ( .D(g29979), .Q(g3060), .CK(CK) );
DFF_X2 U_g3061 ( .D(g30119), .Q(g3061), .CK(CK) );
DFF_X2 U_g3062 ( .D(g30908), .Q(g3062), .CK(CK) );
DFF_X2 U_g3063 ( .D(g30909), .Q(g3063), .CK(CK) );
DFF_X2 U_g3064 ( .D(g30910), .Q(g3064), .CK(CK) );
DFF_X2 U_g3065 ( .D(g30911), .Q(g3065), .CK(CK) );
DFF_X2 U_g3066 ( .D(g30912), .Q(g3066), .CK(CK) );
DFF_X2 U_g3067 ( .D(g30913), .Q(g3067), .CK(CK) );
DFF_X2 U_g3068 ( .D(g30914), .Q(g3068), .CK(CK) );
DFF_X2 U_g3069 ( .D(g30915), .Q(g3069), .CK(CK) );
DFF_X2 U_g3070 ( .D(g30940), .Q(g3070), .CK(CK) );
DFF_X2 U_g3071 ( .D(g30980), .Q(g3071), .CK(CK) );
DFF_X2 U_g3072 ( .D(g30981), .Q(g3072), .CK(CK) );
DFF_X2 U_g3073 ( .D(g30982), .Q(g3073), .CK(CK) );
DFF_X2 U_g3074 ( .D(g30983), .Q(g3074), .CK(CK) );
DFF_X2 U_g3075 ( .D(g30984), .Q(g3075), .CK(CK) );
DFF_X2 U_g3076 ( .D(g30985), .Q(g3076), .CK(CK) );
DFF_X2 U_g3077 ( .D(g30986), .Q(g3077), .CK(CK) );
DFF_X2 U_g3078 ( .D(g30987), .Q(g3078), .CK(CK) );
DFF_X2 U_g2997 ( .D(g30989), .Q(g2997), .CK(CK) );
DFF_X2 U_g2993 ( .D(g26748), .Q(g2993), .CK(CK) );
DFF_X2 U_g2998 ( .D(g27238), .Q(g2998), .CK(CK) );
DFF_X2 U_g3006 ( .D(g25177), .Q(g3006), .CK(CK) );
DFF_X2 U_g3002 ( .D(g26021), .Q(g3002), .CK(CK) );
DFF_X2 U_g3013 ( .D(g26750), .Q(g3013), .CK(CK) );
DFF_X2 U_g3010 ( .D(g27239), .Q(g3010), .CK(CK) );
DFF_X2 U_g3024 ( .D(g27716), .Q(g3024), .CK(CK) );
DFF_X2 U_g3018 ( .D(g24425), .Q(g3018), .CK(CK) );
DFF_X2 U_g3028 ( .D(g25176), .Q(g3028), .CK(CK) );
DFF_X2 U_g3036 ( .D(g26022), .Q(g3036), .CK(CK) );
DFF_X2 U_g3032 ( .D(g26749), .Q(g3032), .CK(CK) );
DFF_X2 U_g3040 ( .D(g16497), .Q(g3040), .CK(CK) );
DFF_X2 U_g2986 ( .D(g3040), .Q(g2986), .CK(CK) );
DFF_X2 U_g2987 ( .D(g16495), .Q(g2987), .CK(CK) );
DFF_X2 U_g48 ( .D(g20595), .Q(g48), .CK(CK) );
DFF_X2 U_g45 ( .D(g20596), .Q(g45), .CK(CK) );
DFF_X2 U_g42 ( .D(g20597), .Q(g42), .CK(CK) );
DFF_X2 U_g39 ( .D(g20598), .Q(g39), .CK(CK) );
DFF_X2 U_g27 ( .D(g20599), .Q(g27), .CK(CK) );
DFF_X2 U_g30 ( .D(g20600), .Q(g30), .CK(CK) );
DFF_X2 U_g33 ( .D(g20601), .Q(g33), .CK(CK) );
DFF_X2 U_g36 ( .D(g20602), .Q(g36), .CK(CK) );
DFF_X2 U_g3083 ( .D(g20603), .Q(g3083), .CK(CK) );
DFF_X2 U_g26 ( .D(g20604), .Q(g26), .CK(CK) );
DFF_X2 U_g2992 ( .D(g21966), .Q(g2992), .CK(CK) );
DFF_X2 U_g23 ( .D(g20605), .Q(g23), .CK(CK) );
DFF_X2 U_g20 ( .D(g20606), .Q(g20), .CK(CK) );
DFF_X2 U_g17 ( .D(g20607), .Q(g17), .CK(CK) );
DFF_X2 U_g11 ( .D(g20608), .Q(g11), .CK(CK) );
DFF_X2 U_g14 ( .D(g20589), .Q(g14), .CK(CK) );
DFF_X2 U_g5 ( .D(g20590), .Q(g5), .CK(CK) );
DFF_X2 U_g8 ( .D(g20591), .Q(g8), .CK(CK) );
DFF_X2 U_g2 ( .D(g20592), .Q(g2), .CK(CK) );
DFF_X2 U_g2990 ( .D(g20593), .Q(g2990), .CK(CK) );
DFF_X2 U_g2991 ( .D(g21964), .Q(g2991), .CK(CK) );
DFF_X2 U_g1 ( .D(g20594), .Q(g1), .CK(CK) );


endmodule

